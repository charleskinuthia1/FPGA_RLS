`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:01:58 04/07/2016 
// Design Name: 
// Module Name:    Gen_K_A 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SignalAKGen(k,a);
	parameter WIDTH = 32;
	
	output [WIDTH*512-1:0] k,a;

	wire [WIDTH*512-1:0] k, a;

	// k values
	assign k[WIDTH*0+:WIDTH]=4860;
	assign k[WIDTH*1+:WIDTH]=-2510;
	assign k[WIDTH*2+:WIDTH]=2937;
	assign k[WIDTH*3+:WIDTH]=11811;
	assign k[WIDTH*4+:WIDTH]=5874;
	assign k[WIDTH*5+:WIDTH]=11249;
	assign k[WIDTH*6+:WIDTH]=-8083;
	assign k[WIDTH*7+:WIDTH]=2661;
	assign k[WIDTH*8+:WIDTH]=-2686;
	assign k[WIDTH*9+:WIDTH]=-2454;
	assign k[WIDTH*10+:WIDTH]=5417;
	assign k[WIDTH*11+:WIDTH]=-6111;
	assign k[WIDTH*12+:WIDTH]=534;
	assign k[WIDTH*13+:WIDTH]=2305;
	assign k[WIDTH*14+:WIDTH]=6680;
	assign k[WIDTH*15+:WIDTH]=6718;
	assign k[WIDTH*16+:WIDTH]=3367;
	assign k[WIDTH*17+:WIDTH]=-3124;
	assign k[WIDTH*18+:WIDTH]=80;
	assign k[WIDTH*19+:WIDTH]=-4410;
	assign k[WIDTH*20+:WIDTH]=-451;
	assign k[WIDTH*21+:WIDTH]=2136;
	assign k[WIDTH*22+:WIDTH]=-5283;
	assign k[WIDTH*23+:WIDTH]=3957;
	assign k[WIDTH*24+:WIDTH]=7174;
	assign k[WIDTH*25+:WIDTH]=-773;
	assign k[WIDTH*26+:WIDTH]=2474;
	assign k[WIDTH*27+:WIDTH]=6067;
	assign k[WIDTH*28+:WIDTH]=-3361;
	assign k[WIDTH*29+:WIDTH]=-3797;
	assign k[WIDTH*30+:WIDTH]=-1259;
	assign k[WIDTH*31+:WIDTH]=7534;
	assign k[WIDTH*32+:WIDTH]=-2217;
	assign k[WIDTH*33+:WIDTH]=3604;
	assign k[WIDTH*34+:WIDTH]=4409;
	assign k[WIDTH*35+:WIDTH]=-1200;
	assign k[WIDTH*36+:WIDTH]=-7864;
	assign k[WIDTH*37+:WIDTH]=5310;
	assign k[WIDTH*38+:WIDTH]=-8018;
	assign k[WIDTH*39+:WIDTH]=-11380;
	assign k[WIDTH*40+:WIDTH]=470;
	assign k[WIDTH*41+:WIDTH]=-13707;
	assign k[WIDTH*42+:WIDTH]=-8941;
	assign k[WIDTH*43+:WIDTH]=-6606;
	assign k[WIDTH*44+:WIDTH]=8630;
	assign k[WIDTH*45+:WIDTH]=240;
	assign k[WIDTH*46+:WIDTH]=-5961;
	assign k[WIDTH*47+:WIDTH]=4808;
	assign k[WIDTH*48+:WIDTH]=2517;
	assign k[WIDTH*49+:WIDTH]=9935;
	assign k[WIDTH*50+:WIDTH]=4806;
	assign k[WIDTH*51+:WIDTH]=-7644;
	assign k[WIDTH*52+:WIDTH]=4042;
	assign k[WIDTH*53+:WIDTH]=-3379;
	assign k[WIDTH*54+:WIDTH]=6777;
	assign k[WIDTH*55+:WIDTH]=-2778;
	assign k[WIDTH*56+:WIDTH]=3008;
	assign k[WIDTH*57+:WIDTH]=4498;
	assign k[WIDTH*58+:WIDTH]=5755;
	assign k[WIDTH*59+:WIDTH]=9950;
	assign k[WIDTH*60+:WIDTH]=10057;
	assign k[WIDTH*61+:WIDTH]=2035;
	assign k[WIDTH*62+:WIDTH]=2307;
	assign k[WIDTH*63+:WIDTH]=854;
	assign k[WIDTH*64+:WIDTH]=391;
	assign k[WIDTH*65+:WIDTH]=9270;
	assign k[WIDTH*66+:WIDTH]=-8833;
	assign k[WIDTH*67+:WIDTH]=3370;
	assign k[WIDTH*68+:WIDTH]=-8735;
	assign k[WIDTH*69+:WIDTH]=8548;
	assign k[WIDTH*70+:WIDTH]=7508;
	assign k[WIDTH*71+:WIDTH]=-6797;
	assign k[WIDTH*72+:WIDTH]=3407;
	assign k[WIDTH*73+:WIDTH]=-2707;
	assign k[WIDTH*74+:WIDTH]=1819;
	assign k[WIDTH*75+:WIDTH]=5494;
	assign k[WIDTH*76+:WIDTH]=2931;
	assign k[WIDTH*77+:WIDTH]=1387;
	assign k[WIDTH*78+:WIDTH]=4175;
	assign k[WIDTH*79+:WIDTH]=1478;
	assign k[WIDTH*80+:WIDTH]=-9725;
	assign k[WIDTH*81+:WIDTH]=3170;
	assign k[WIDTH*82+:WIDTH]=4578;
	assign k[WIDTH*83+:WIDTH]=1687;
	assign k[WIDTH*84+:WIDTH]=-6325;
	assign k[WIDTH*85+:WIDTH]=-1257;
	assign k[WIDTH*86+:WIDTH]=-7061;
	assign k[WIDTH*87+:WIDTH]=49;
	assign k[WIDTH*88+:WIDTH]=3271;
	assign k[WIDTH*89+:WIDTH]=10730;
	assign k[WIDTH*90+:WIDTH]=-2923;
	assign k[WIDTH*91+:WIDTH]=2957;
	assign k[WIDTH*92+:WIDTH]=3629;
	assign k[WIDTH*93+:WIDTH]=4820;
	assign k[WIDTH*94+:WIDTH]=4380;
	assign k[WIDTH*95+:WIDTH]=2870;
	assign k[WIDTH*96+:WIDTH]=4380;
	assign k[WIDTH*97+:WIDTH]=9269;
	assign k[WIDTH*98+:WIDTH]=4322;
	assign k[WIDTH*99+:WIDTH]=3484;
	assign k[WIDTH*100+:WIDTH]=-2240;
	assign k[WIDTH*101+:WIDTH]=-2964;
	assign k[WIDTH*102+:WIDTH]=-6268;
	assign k[WIDTH*103+:WIDTH]=2973;
	assign k[WIDTH*104+:WIDTH]=-3613;
	assign k[WIDTH*105+:WIDTH]=706;
	assign k[WIDTH*106+:WIDTH]=10616;
	assign k[WIDTH*107+:WIDTH]=890;
	assign k[WIDTH*108+:WIDTH]=-8609;
	assign k[WIDTH*109+:WIDTH]=1057;
	assign k[WIDTH*110+:WIDTH]=-1824;
	assign k[WIDTH*111+:WIDTH]=-5989;
	assign k[WIDTH*112+:WIDTH]=-1396;
	assign k[WIDTH*113+:WIDTH]=-2465;
	assign k[WIDTH*114+:WIDTH]=-2383;
	assign k[WIDTH*115+:WIDTH]=-4501;
	assign k[WIDTH*116+:WIDTH]=8873;
	assign k[WIDTH*117+:WIDTH]=7071;
	assign k[WIDTH*118+:WIDTH]=-7810;
	assign k[WIDTH*119+:WIDTH]=6144;
	assign k[WIDTH*120+:WIDTH]=-653;
	assign k[WIDTH*121+:WIDTH]=-1546;
	assign k[WIDTH*122+:WIDTH]=1525;
	assign k[WIDTH*123+:WIDTH]=-5418;
	assign k[WIDTH*124+:WIDTH]=222;
	assign k[WIDTH*125+:WIDTH]=6143;
	assign k[WIDTH*126+:WIDTH]=-489;
	assign k[WIDTH*127+:WIDTH]=-14939;
	assign k[WIDTH*128+:WIDTH]=3479;
	assign k[WIDTH*129+:WIDTH]=4596;
	assign k[WIDTH*130+:WIDTH]=9629;
	assign k[WIDTH*131+:WIDTH]=-3167;
	assign k[WIDTH*132+:WIDTH]=-7267;
	assign k[WIDTH*133+:WIDTH]=4456;
	assign k[WIDTH*134+:WIDTH]=8610;
	assign k[WIDTH*135+:WIDTH]=2197;
	assign k[WIDTH*136+:WIDTH]=3792;
	assign k[WIDTH*137+:WIDTH]=-2256;
	assign k[WIDTH*138+:WIDTH]=-2532;
	assign k[WIDTH*139+:WIDTH]=-1742;
	assign k[WIDTH*140+:WIDTH]=-3682;
	assign k[WIDTH*141+:WIDTH]=-4482;
	assign k[WIDTH*142+:WIDTH]=5663;
	assign k[WIDTH*143+:WIDTH]=-4335;
	assign k[WIDTH*144+:WIDTH]=-540;
	assign k[WIDTH*145+:WIDTH]=-3756;
	assign k[WIDTH*146+:WIDTH]=2046;
	assign k[WIDTH*147+:WIDTH]=18069;
	assign k[WIDTH*148+:WIDTH]=1153;
	assign k[WIDTH*149+:WIDTH]=7639;
	assign k[WIDTH*150+:WIDTH]=10207;
	assign k[WIDTH*151+:WIDTH]=9745;
	assign k[WIDTH*152+:WIDTH]=13504;
	assign k[WIDTH*153+:WIDTH]=13302;
	assign k[WIDTH*154+:WIDTH]=8890;
	assign k[WIDTH*155+:WIDTH]=641;
	assign k[WIDTH*156+:WIDTH]=1886;
	assign k[WIDTH*157+:WIDTH]=11525;
	assign k[WIDTH*158+:WIDTH]=-32143;
	assign k[WIDTH*159+:WIDTH]=-1904;
	assign k[WIDTH*160+:WIDTH]=12982;
	assign k[WIDTH*161+:WIDTH]=-1425;
	assign k[WIDTH*162+:WIDTH]=8157;
	assign k[WIDTH*163+:WIDTH]=8408;
	assign k[WIDTH*164+:WIDTH]=-10135;
	assign k[WIDTH*165+:WIDTH]=-3539;
	assign k[WIDTH*166+:WIDTH]=1941;
	assign k[WIDTH*167+:WIDTH]=10464;
	assign k[WIDTH*168+:WIDTH]=-5730;
	assign k[WIDTH*169+:WIDTH]=-21613;
	assign k[WIDTH*170+:WIDTH]=-5476;
	assign k[WIDTH*171+:WIDTH]=11362;
	assign k[WIDTH*172+:WIDTH]=3971;
	assign k[WIDTH*173+:WIDTH]=1122;
	assign k[WIDTH*174+:WIDTH]=1331;
	assign k[WIDTH*175+:WIDTH]=-4831;
	assign k[WIDTH*176+:WIDTH]=-2764;
	assign k[WIDTH*177+:WIDTH]=461;
	assign k[WIDTH*178+:WIDTH]=-3986;
	assign k[WIDTH*179+:WIDTH]=5446;
	assign k[WIDTH*180+:WIDTH]=3689;
	assign k[WIDTH*181+:WIDTH]=-10270;
	assign k[WIDTH*182+:WIDTH]=2773;
	assign k[WIDTH*183+:WIDTH]=10203;
	assign k[WIDTH*184+:WIDTH]=8453;
	assign k[WIDTH*185+:WIDTH]=-3026;
	assign k[WIDTH*186+:WIDTH]=-850;
	assign k[WIDTH*187+:WIDTH]=-6965;
	assign k[WIDTH*188+:WIDTH]=5021;
	assign k[WIDTH*189+:WIDTH]=464;
	assign k[WIDTH*190+:WIDTH]=719;
	assign k[WIDTH*191+:WIDTH]=1525;
	assign k[WIDTH*192+:WIDTH]=-10206;
	assign k[WIDTH*193+:WIDTH]=14661;
	assign k[WIDTH*194+:WIDTH]=1614;
	assign k[WIDTH*195+:WIDTH]=-2566;
	assign k[WIDTH*196+:WIDTH]=11047;
	assign k[WIDTH*197+:WIDTH]=9649;
	assign k[WIDTH*198+:WIDTH]=-6472;
	assign k[WIDTH*199+:WIDTH]=-10889;
	assign k[WIDTH*200+:WIDTH]=-5485;
	assign k[WIDTH*201+:WIDTH]=12055;
	assign k[WIDTH*202+:WIDTH]=-13303;
	assign k[WIDTH*203+:WIDTH]=13841;
	assign k[WIDTH*204+:WIDTH]=-6856;
	assign k[WIDTH*205+:WIDTH]=-15182;
	assign k[WIDTH*206+:WIDTH]=-9135;
	assign k[WIDTH*207+:WIDTH]=3445;
	assign k[WIDTH*208+:WIDTH]=-4940;
	assign k[WIDTH*209+:WIDTH]=-3914;
	assign k[WIDTH*210+:WIDTH]=14623;
	assign k[WIDTH*211+:WIDTH]=-9353;
	assign k[WIDTH*212+:WIDTH]=3085;
	assign k[WIDTH*213+:WIDTH]=4785;
	assign k[WIDTH*214+:WIDTH]=1874;
	assign k[WIDTH*215+:WIDTH]=-2942;
	assign k[WIDTH*216+:WIDTH]=-4558;
	assign k[WIDTH*217+:WIDTH]=-9473;
	assign k[WIDTH*218+:WIDTH]=-1071;
	assign k[WIDTH*219+:WIDTH]=-3393;
	assign k[WIDTH*220+:WIDTH]=-9416;
	assign k[WIDTH*221+:WIDTH]=24377;
	assign k[WIDTH*222+:WIDTH]=-70;
	assign k[WIDTH*223+:WIDTH]=10138;
	assign k[WIDTH*224+:WIDTH]=-12337;
	assign k[WIDTH*225+:WIDTH]=1255;
	assign k[WIDTH*226+:WIDTH]=9611;
	assign k[WIDTH*227+:WIDTH]=-1494;
	assign k[WIDTH*228+:WIDTH]=2701;
	assign k[WIDTH*229+:WIDTH]=4846;
	assign k[WIDTH*230+:WIDTH]=4041;
	assign k[WIDTH*231+:WIDTH]=8331;
	assign k[WIDTH*232+:WIDTH]=-4634;
	assign k[WIDTH*233+:WIDTH]=-12907;
	assign k[WIDTH*234+:WIDTH]=3311;
	assign k[WIDTH*235+:WIDTH]=1502;
	assign k[WIDTH*236+:WIDTH]=-1301;
	assign k[WIDTH*237+:WIDTH]=5553;
	assign k[WIDTH*238+:WIDTH]=-11722;
	assign k[WIDTH*239+:WIDTH]=6102;
	assign k[WIDTH*240+:WIDTH]=8200;
	assign k[WIDTH*241+:WIDTH]=4566;
	assign k[WIDTH*242+:WIDTH]=-118;
	assign k[WIDTH*243+:WIDTH]=20736;
	assign k[WIDTH*244+:WIDTH]=-2622;
	assign k[WIDTH*245+:WIDTH]=-10161;
	assign k[WIDTH*246+:WIDTH]=-945;
	assign k[WIDTH*247+:WIDTH]=-13349;
	assign k[WIDTH*248+:WIDTH]=12947;
	assign k[WIDTH*249+:WIDTH]=-1324;
	assign k[WIDTH*250+:WIDTH]=-11885;
	assign k[WIDTH*251+:WIDTH]=15879;
	assign k[WIDTH*252+:WIDTH]=-12009;
	assign k[WIDTH*253+:WIDTH]=2947;
	assign k[WIDTH*254+:WIDTH]=11121;
	assign k[WIDTH*255+:WIDTH]=-9672;
	assign k[WIDTH*256+:WIDTH]=-28683;
	assign k[WIDTH*257+:WIDTH]=-9165;
	assign k[WIDTH*258+:WIDTH]=8093;
	assign k[WIDTH*259+:WIDTH]=-9013;
	assign k[WIDTH*260+:WIDTH]=7862;
	assign k[WIDTH*261+:WIDTH]=3483;
	assign k[WIDTH*262+:WIDTH]=1493;
	assign k[WIDTH*263+:WIDTH]=-11303;
	assign k[WIDTH*264+:WIDTH]=776;
	assign k[WIDTH*265+:WIDTH]=-10140;
	assign k[WIDTH*266+:WIDTH]=18984;
	assign k[WIDTH*267+:WIDTH]=2359;
	assign k[WIDTH*268+:WIDTH]=472;
	assign k[WIDTH*269+:WIDTH]=-9388;
	assign k[WIDTH*270+:WIDTH]=-7404;
	assign k[WIDTH*271+:WIDTH]=5463;
	assign k[WIDTH*272+:WIDTH]=-250;
	assign k[WIDTH*273+:WIDTH]=-7744;
	assign k[WIDTH*274+:WIDTH]=-2744;
	assign k[WIDTH*275+:WIDTH]=921;
	assign k[WIDTH*276+:WIDTH]=-8465;
	assign k[WIDTH*277+:WIDTH]=-3671;
	assign k[WIDTH*278+:WIDTH]=4415;
	assign k[WIDTH*279+:WIDTH]=-2616;
	assign k[WIDTH*280+:WIDTH]=8284;
	assign k[WIDTH*281+:WIDTH]=-2499;
	assign k[WIDTH*282+:WIDTH]=9179;
	assign k[WIDTH*283+:WIDTH]=-4281;
	assign k[WIDTH*284+:WIDTH]=-2164;
	assign k[WIDTH*285+:WIDTH]=7803;
	assign k[WIDTH*286+:WIDTH]=12146;
	assign k[WIDTH*287+:WIDTH]=-6306;
	assign k[WIDTH*288+:WIDTH]=-7361;
	assign k[WIDTH*289+:WIDTH]=-8474;
	assign k[WIDTH*290+:WIDTH]=608;
	assign k[WIDTH*291+:WIDTH]=-10866;
	assign k[WIDTH*292+:WIDTH]=-8360;
	assign k[WIDTH*293+:WIDTH]=2269;
	assign k[WIDTH*294+:WIDTH]=3628;
	assign k[WIDTH*295+:WIDTH]=2799;
	assign k[WIDTH*296+:WIDTH]=866;
	assign k[WIDTH*297+:WIDTH]=-1808;
	assign k[WIDTH*298+:WIDTH]=20702;
	assign k[WIDTH*299+:WIDTH]=-13435;
	assign k[WIDTH*300+:WIDTH]=5424;
	assign k[WIDTH*301+:WIDTH]=748;
	assign k[WIDTH*302+:WIDTH]=1174;
	assign k[WIDTH*303+:WIDTH]=3128;
	assign k[WIDTH*304+:WIDTH]=13420;
	assign k[WIDTH*305+:WIDTH]=2715;
	assign k[WIDTH*306+:WIDTH]=-2500;
	assign k[WIDTH*307+:WIDTH]=593;
	assign k[WIDTH*308+:WIDTH]=-2818;
	assign k[WIDTH*309+:WIDTH]=-1600;
	assign k[WIDTH*310+:WIDTH]=-2076;
	assign k[WIDTH*311+:WIDTH]=7831;
	assign k[WIDTH*312+:WIDTH]=-2265;
	assign k[WIDTH*313+:WIDTH]=1486;
	assign k[WIDTH*314+:WIDTH]=-11622;
	assign k[WIDTH*315+:WIDTH]=-6864;
	assign k[WIDTH*316+:WIDTH]=-2984;
	assign k[WIDTH*317+:WIDTH]=9580;
	assign k[WIDTH*318+:WIDTH]=9641;
	assign k[WIDTH*319+:WIDTH]=-221;
	assign k[WIDTH*320+:WIDTH]=5563;
	assign k[WIDTH*321+:WIDTH]=7065;
	assign k[WIDTH*322+:WIDTH]=-1160;
	assign k[WIDTH*323+:WIDTH]=1956;
	assign k[WIDTH*324+:WIDTH]=-578;
	assign k[WIDTH*325+:WIDTH]=-1433;
	assign k[WIDTH*326+:WIDTH]=-592;
	assign k[WIDTH*327+:WIDTH]=4966;
	assign k[WIDTH*328+:WIDTH]=-706;
	assign k[WIDTH*329+:WIDTH]=1500;
	assign k[WIDTH*330+:WIDTH]=-12113;
	assign k[WIDTH*331+:WIDTH]=-316;
	assign k[WIDTH*332+:WIDTH]=-4252;
	assign k[WIDTH*333+:WIDTH]=4653;
	assign k[WIDTH*334+:WIDTH]=5716;
	assign k[WIDTH*335+:WIDTH]=1761;
	assign k[WIDTH*336+:WIDTH]=-6602;
	assign k[WIDTH*337+:WIDTH]=3612;
	assign k[WIDTH*338+:WIDTH]=3517;
	assign k[WIDTH*339+:WIDTH]=-4143;
	assign k[WIDTH*340+:WIDTH]=-2382;
	assign k[WIDTH*341+:WIDTH]=626;
	assign k[WIDTH*342+:WIDTH]=569;
	assign k[WIDTH*343+:WIDTH]=9188;
	assign k[WIDTH*344+:WIDTH]=-5623;
	assign k[WIDTH*345+:WIDTH]=-4776;
	assign k[WIDTH*346+:WIDTH]=9880;
	assign k[WIDTH*347+:WIDTH]=-4269;
	assign k[WIDTH*348+:WIDTH]=2672;
	assign k[WIDTH*349+:WIDTH]=-3146;
	assign k[WIDTH*350+:WIDTH]=-5926;
	assign k[WIDTH*351+:WIDTH]=4092;
	assign k[WIDTH*352+:WIDTH]=7264;
	assign k[WIDTH*353+:WIDTH]=-3637;
	assign k[WIDTH*354+:WIDTH]=-1073;
	assign k[WIDTH*355+:WIDTH]=-4046;
	assign k[WIDTH*356+:WIDTH]=-6770;
	assign k[WIDTH*357+:WIDTH]=-3562;
	assign k[WIDTH*358+:WIDTH]=3834;
	assign k[WIDTH*359+:WIDTH]=3298;
	assign k[WIDTH*360+:WIDTH]=10;
	assign k[WIDTH*361+:WIDTH]=1053;
	assign k[WIDTH*362+:WIDTH]=3273;
	assign k[WIDTH*363+:WIDTH]=-5952;
	assign k[WIDTH*364+:WIDTH]=4393;
	assign k[WIDTH*365+:WIDTH]=8429;
	assign k[WIDTH*366+:WIDTH]=-1897;
	assign k[WIDTH*367+:WIDTH]=2345;
	assign k[WIDTH*368+:WIDTH]=1956;
	assign k[WIDTH*369+:WIDTH]=3933;
	assign k[WIDTH*370+:WIDTH]=1450;
	assign k[WIDTH*371+:WIDTH]=-494;
	assign k[WIDTH*372+:WIDTH]=1936;
	assign k[WIDTH*373+:WIDTH]=-3669;
	assign k[WIDTH*374+:WIDTH]=631;
	assign k[WIDTH*375+:WIDTH]=-5458;
	assign k[WIDTH*376+:WIDTH]=501;
	assign k[WIDTH*377+:WIDTH]=-557;
	assign k[WIDTH*378+:WIDTH]=-5615;
	assign k[WIDTH*379+:WIDTH]=-1649;
	assign k[WIDTH*380+:WIDTH]=-8132;
	assign k[WIDTH*381+:WIDTH]=5993;
	assign k[WIDTH*382+:WIDTH]=616;
	assign k[WIDTH*383+:WIDTH]=2753;
	assign k[WIDTH*384+:WIDTH]=-2209;
	assign k[WIDTH*385+:WIDTH]=2411;
	assign k[WIDTH*386+:WIDTH]=5654;
	assign k[WIDTH*387+:WIDTH]=7655;
	assign k[WIDTH*388+:WIDTH]=6608;
	assign k[WIDTH*389+:WIDTH]=1612;
	assign k[WIDTH*390+:WIDTH]=869;
	assign k[WIDTH*391+:WIDTH]=719;
	assign k[WIDTH*392+:WIDTH]=1573;
	assign k[WIDTH*393+:WIDTH]=-1409;
	assign k[WIDTH*394+:WIDTH]=-1991;
	assign k[WIDTH*395+:WIDTH]=8501;
	assign k[WIDTH*396+:WIDTH]=-758;
	assign k[WIDTH*397+:WIDTH]=930;
	assign k[WIDTH*398+:WIDTH]=-2899;
	assign k[WIDTH*399+:WIDTH]=-3430;
	assign k[WIDTH*400+:WIDTH]=-3430;
	assign k[WIDTH*401+:WIDTH]=-888;
	assign k[WIDTH*402+:WIDTH]=1358;
	assign k[WIDTH*403+:WIDTH]=1484;
	assign k[WIDTH*404+:WIDTH]=1605;
	assign k[WIDTH*405+:WIDTH]=-4088;
	assign k[WIDTH*406+:WIDTH]=-951;
	assign k[WIDTH*407+:WIDTH]=248;
	assign k[WIDTH*408+:WIDTH]=-3655;
	assign k[WIDTH*409+:WIDTH]=-3698;
	assign k[WIDTH*410+:WIDTH]=5331;
	assign k[WIDTH*411+:WIDTH]=3707;
	assign k[WIDTH*412+:WIDTH]=4045;
	assign k[WIDTH*413+:WIDTH]=387;
	assign k[WIDTH*414+:WIDTH]=-798;
	assign k[WIDTH*415+:WIDTH]=1003;
	assign k[WIDTH*416+:WIDTH]=3819;
	assign k[WIDTH*417+:WIDTH]=-3151;
	assign k[WIDTH*418+:WIDTH]=1033;
	assign k[WIDTH*419+:WIDTH]=1555;
	assign k[WIDTH*420+:WIDTH]=710;
	assign k[WIDTH*421+:WIDTH]=785;
	assign k[WIDTH*422+:WIDTH]=3982;
	assign k[WIDTH*423+:WIDTH]=-6420;
	assign k[WIDTH*424+:WIDTH]=1542;
	assign k[WIDTH*425+:WIDTH]=6928;
	assign k[WIDTH*426+:WIDTH]=-1298;
	assign k[WIDTH*427+:WIDTH]=1971;
	assign k[WIDTH*428+:WIDTH]=-1458;
	assign k[WIDTH*429+:WIDTH]=3516;
	assign k[WIDTH*430+:WIDTH]=1097;
	assign k[WIDTH*431+:WIDTH]=2177;
	assign k[WIDTH*432+:WIDTH]=-1931;
	assign k[WIDTH*433+:WIDTH]=-1640;
	assign k[WIDTH*434+:WIDTH]=-150;
	assign k[WIDTH*435+:WIDTH]=-165;
	assign k[WIDTH*436+:WIDTH]=-3182;
	assign k[WIDTH*437+:WIDTH]=5908;
	assign k[WIDTH*438+:WIDTH]=2105;
	assign k[WIDTH*439+:WIDTH]=4850;
	assign k[WIDTH*440+:WIDTH]=-6456;
	assign k[WIDTH*441+:WIDTH]=4303;
	assign k[WIDTH*442+:WIDTH]=674;
	assign k[WIDTH*443+:WIDTH]=-1010;
	assign k[WIDTH*444+:WIDTH]=-1312;
	assign k[WIDTH*445+:WIDTH]=1424;
	assign k[WIDTH*446+:WIDTH]=-1661;
	assign k[WIDTH*447+:WIDTH]=1111;
	assign k[WIDTH*448+:WIDTH]=8921;
	assign k[WIDTH*449+:WIDTH]=-2798;
	assign k[WIDTH*450+:WIDTH]=2655;
	assign k[WIDTH*451+:WIDTH]=2231;
	assign k[WIDTH*452+:WIDTH]=-1613;
	assign k[WIDTH*453+:WIDTH]=1544;
	assign k[WIDTH*454+:WIDTH]=-2005;
	assign k[WIDTH*455+:WIDTH]=-3227;
	assign k[WIDTH*456+:WIDTH]=1056;
	assign k[WIDTH*457+:WIDTH]=6871;
	assign k[WIDTH*458+:WIDTH]=-546;
	assign k[WIDTH*459+:WIDTH]=1529;
	assign k[WIDTH*460+:WIDTH]=1962;
	assign k[WIDTH*461+:WIDTH]=-2070;
	assign k[WIDTH*462+:WIDTH]=-1369;
	assign k[WIDTH*463+:WIDTH]=1287;
	assign k[WIDTH*464+:WIDTH]=-4011;
	assign k[WIDTH*465+:WIDTH]=1318;
	assign k[WIDTH*466+:WIDTH]=-4769;
	assign k[WIDTH*467+:WIDTH]=-4115;
	assign k[WIDTH*468+:WIDTH]=909;
	assign k[WIDTH*469+:WIDTH]=2157;
	assign k[WIDTH*470+:WIDTH]=-2570;
	assign k[WIDTH*471+:WIDTH]=2442;
	assign k[WIDTH*472+:WIDTH]=-3020;
	assign k[WIDTH*473+:WIDTH]=234;
	assign k[WIDTH*474+:WIDTH]=-4662;
	assign k[WIDTH*475+:WIDTH]=-1789;
	assign k[WIDTH*476+:WIDTH]=-2173;
	assign k[WIDTH*477+:WIDTH]=-45;
	assign k[WIDTH*478+:WIDTH]=110;
	assign k[WIDTH*479+:WIDTH]=1885;
	assign k[WIDTH*480+:WIDTH]=7827;
	assign k[WIDTH*481+:WIDTH]=-1406;
	assign k[WIDTH*482+:WIDTH]=-71;
	assign k[WIDTH*483+:WIDTH]=-3629;
	assign k[WIDTH*484+:WIDTH]=-2932;
	assign k[WIDTH*485+:WIDTH]=1913;
	assign k[WIDTH*486+:WIDTH]=-869;
	assign k[WIDTH*487+:WIDTH]=-591;
	assign k[WIDTH*488+:WIDTH]=-3280;
	assign k[WIDTH*489+:WIDTH]=6705;
	assign k[WIDTH*490+:WIDTH]=-2215;
	assign k[WIDTH*491+:WIDTH]=-2220;
	assign k[WIDTH*492+:WIDTH]=798;
	assign k[WIDTH*493+:WIDTH]=2114;
	assign k[WIDTH*494+:WIDTH]=-4316;
	assign k[WIDTH*495+:WIDTH]=2654;
	assign k[WIDTH*496+:WIDTH]=-7212;
	assign k[WIDTH*497+:WIDTH]=3207;
	assign k[WIDTH*498+:WIDTH]=-1341;
	assign k[WIDTH*499+:WIDTH]=-4232;
	assign k[WIDTH*500+:WIDTH]=311;
	assign k[WIDTH*501+:WIDTH]=-208;
	assign k[WIDTH*502+:WIDTH]=3009;
	assign k[WIDTH*503+:WIDTH]=1107;
	assign k[WIDTH*504+:WIDTH]=-3105;
	assign k[WIDTH*505+:WIDTH]=-4116;
	assign k[WIDTH*506+:WIDTH]=4059;
	assign k[WIDTH*507+:WIDTH]=-3043;
	assign k[WIDTH*508+:WIDTH]=-3039;
	assign k[WIDTH*509+:WIDTH]=460;
	assign k[WIDTH*510+:WIDTH]=-555;
	assign k[WIDTH*511+:WIDTH]=5778;

	
	// a values
		assign a[WIDTH*0+:WIDTH]=32998;
	assign a[WIDTH*1+:WIDTH]=-2228;
	assign a[WIDTH*2+:WIDTH]=58444;
	assign a[WIDTH*3+:WIDTH]=98690;
	assign a[WIDTH*4+:WIDTH]=76307;
	assign a[WIDTH*5+:WIDTH]=80562;
	assign a[WIDTH*6+:WIDTH]=-18563;
	assign a[WIDTH*7+:WIDTH]=581;
	assign a[WIDTH*8+:WIDTH]=-13736;
	assign a[WIDTH*9+:WIDTH]=5512;
	assign a[WIDTH*10+:WIDTH]=38628;
	assign a[WIDTH*11+:WIDTH]=-31227;
	assign a[WIDTH*12+:WIDTH]=41823;
	assign a[WIDTH*13+:WIDTH]=-20255;
	assign a[WIDTH*14+:WIDTH]=73403;
	assign a[WIDTH*15+:WIDTH]=56904;
	assign a[WIDTH*16+:WIDTH]=65170;
	assign a[WIDTH*17+:WIDTH]=-24703;
	assign a[WIDTH*18+:WIDTH]=-21575;
	assign a[WIDTH*19+:WIDTH]=-76494;
	assign a[WIDTH*20+:WIDTH]=222;
	assign a[WIDTH*21+:WIDTH]=60511;
	assign a[WIDTH*22+:WIDTH]=-108328;
	assign a[WIDTH*23+:WIDTH]=66683;
	assign a[WIDTH*24+:WIDTH]=158028;
	assign a[WIDTH*25+:WIDTH]=-32210;
	assign a[WIDTH*26+:WIDTH]=29184;
	assign a[WIDTH*27+:WIDTH]=71992;
	assign a[WIDTH*28+:WIDTH]=-51808;
	assign a[WIDTH*29+:WIDTH]=-29232;
	assign a[WIDTH*30+:WIDTH]=-159;
	assign a[WIDTH*31+:WIDTH]=98005;
	assign a[WIDTH*32+:WIDTH]=-2205;
	assign a[WIDTH*33+:WIDTH]=59338;
	assign a[WIDTH*34+:WIDTH]=43904;
	assign a[WIDTH*35+:WIDTH]=19599;
	assign a[WIDTH*36+:WIDTH]=-28975;
	assign a[WIDTH*37+:WIDTH]=-42405;
	assign a[WIDTH*38+:WIDTH]=-13724;
	assign a[WIDTH*39+:WIDTH]=-115943;
	assign a[WIDTH*40+:WIDTH]=-28861;
	assign a[WIDTH*41+:WIDTH]=-34672;
	assign a[WIDTH*42+:WIDTH]=-42752;
	assign a[WIDTH*43+:WIDTH]=-108312;
	assign a[WIDTH*44+:WIDTH]=83315;
	assign a[WIDTH*45+:WIDTH]=12036;
	assign a[WIDTH*46+:WIDTH]=-71447;
	assign a[WIDTH*47+:WIDTH]=-52456;
	assign a[WIDTH*48+:WIDTH]=19269;
	assign a[WIDTH*49+:WIDTH]=19019;
	assign a[WIDTH*50+:WIDTH]=-3225;
	assign a[WIDTH*51+:WIDTH]=-107463;
	assign a[WIDTH*52+:WIDTH]=60436;
	assign a[WIDTH*53+:WIDTH]=-67216;
	assign a[WIDTH*54+:WIDTH]=83027;
	assign a[WIDTH*55+:WIDTH]=41945;
	assign a[WIDTH*56+:WIDTH]=6833;
	assign a[WIDTH*57+:WIDTH]=51787;
	assign a[WIDTH*58+:WIDTH]=42570;
	assign a[WIDTH*59+:WIDTH]=137255;
	assign a[WIDTH*60+:WIDTH]=33832;
	assign a[WIDTH*61+:WIDTH]=44291;
	assign a[WIDTH*62+:WIDTH]=20426;
	assign a[WIDTH*63+:WIDTH]=-27230;
	assign a[WIDTH*64+:WIDTH]=25252;
	assign a[WIDTH*65+:WIDTH]=149406;
	assign a[WIDTH*66+:WIDTH]=-52591;
	assign a[WIDTH*67+:WIDTH]=27853;
	assign a[WIDTH*68+:WIDTH]=21147;
	assign a[WIDTH*69+:WIDTH]=103586;
	assign a[WIDTH*70+:WIDTH]=10220;
	assign a[WIDTH*71+:WIDTH]=-60218;
	assign a[WIDTH*72+:WIDTH]=48379;
	assign a[WIDTH*73+:WIDTH]=-62560;
	assign a[WIDTH*74+:WIDTH]=63460;
	assign a[WIDTH*75+:WIDTH]=8597;
	assign a[WIDTH*76+:WIDTH]=117153;
	assign a[WIDTH*77+:WIDTH]=55167;
	assign a[WIDTH*78+:WIDTH]=42114;
	assign a[WIDTH*79+:WIDTH]=35486;
	assign a[WIDTH*80+:WIDTH]=-98215;
	assign a[WIDTH*81+:WIDTH]=22228;
	assign a[WIDTH*82+:WIDTH]=79910;
	assign a[WIDTH*83+:WIDTH]=16861;
	assign a[WIDTH*84+:WIDTH]=-104211;
	assign a[WIDTH*85+:WIDTH]=-17896;
	assign a[WIDTH*86+:WIDTH]=-90004;
	assign a[WIDTH*87+:WIDTH]=10200;
	assign a[WIDTH*88+:WIDTH]=5876;
	assign a[WIDTH*89+:WIDTH]=68037;
	assign a[WIDTH*90+:WIDTH]=-34580;
	assign a[WIDTH*91+:WIDTH]=12790;
	assign a[WIDTH*92+:WIDTH]=103360;
	assign a[WIDTH*93+:WIDTH]=49540;
	assign a[WIDTH*94+:WIDTH]=27022;
	assign a[WIDTH*95+:WIDTH]=-25709;
	assign a[WIDTH*96+:WIDTH]=60023;
	assign a[WIDTH*97+:WIDTH]=10184;
	assign a[WIDTH*98+:WIDTH]=81645;
	assign a[WIDTH*99+:WIDTH]=-36580;
	assign a[WIDTH*100+:WIDTH]=43007;
	assign a[WIDTH*101+:WIDTH]=-126347;
	assign a[WIDTH*102+:WIDTH]=-62647;
	assign a[WIDTH*103+:WIDTH]=100107;
	assign a[WIDTH*104+:WIDTH]=-25766;
	assign a[WIDTH*105+:WIDTH]=66527;
	assign a[WIDTH*106+:WIDTH]=122564;
	assign a[WIDTH*107+:WIDTH]=47807;
	assign a[WIDTH*108+:WIDTH]=-149224;
	assign a[WIDTH*109+:WIDTH]=-38720;
	assign a[WIDTH*110+:WIDTH]=-6813;
	assign a[WIDTH*111+:WIDTH]=1316;
	assign a[WIDTH*112+:WIDTH]=-2590;
	assign a[WIDTH*113+:WIDTH]=1036;
	assign a[WIDTH*114+:WIDTH]=23462;
	assign a[WIDTH*115+:WIDTH]=-71126;
	assign a[WIDTH*116+:WIDTH]=66430;
	assign a[WIDTH*117+:WIDTH]=-40751;
	assign a[WIDTH*118+:WIDTH]=-61594;
	assign a[WIDTH*119+:WIDTH]=44507;
	assign a[WIDTH*120+:WIDTH]=-2763;
	assign a[WIDTH*121+:WIDTH]=-3404;
	assign a[WIDTH*122+:WIDTH]=13161;
	assign a[WIDTH*123+:WIDTH]=-9215;
	assign a[WIDTH*124+:WIDTH]=-46935;
	assign a[WIDTH*125+:WIDTH]=22038;
	assign a[WIDTH*126+:WIDTH]=-35018;
	assign a[WIDTH*127+:WIDTH]=-183233;
	assign a[WIDTH*128+:WIDTH]=17453;
	assign a[WIDTH*129+:WIDTH]=27242;
	assign a[WIDTH*130+:WIDTH]=121280;
	assign a[WIDTH*131+:WIDTH]=-83668;
	assign a[WIDTH*132+:WIDTH]=9502;
	assign a[WIDTH*133+:WIDTH]=-15173;
	assign a[WIDTH*134+:WIDTH]=174273;
	assign a[WIDTH*135+:WIDTH]=17434;
	assign a[WIDTH*136+:WIDTH]=37236;
	assign a[WIDTH*137+:WIDTH]=31413;
	assign a[WIDTH*138+:WIDTH]=-34252;
	assign a[WIDTH*139+:WIDTH]=-44343;
	assign a[WIDTH*140+:WIDTH]=-47690;
	assign a[WIDTH*141+:WIDTH]=-67823;
	assign a[WIDTH*142+:WIDTH]=12583;
	assign a[WIDTH*143+:WIDTH]=-110694;
	assign a[WIDTH*144+:WIDTH]=45522;
	assign a[WIDTH*145+:WIDTH]=-75239;
	assign a[WIDTH*146+:WIDTH]=1341;
	assign a[WIDTH*147+:WIDTH]=4663;
	assign a[WIDTH*148+:WIDTH]=-25;
	assign a[WIDTH*149+:WIDTH]=29806;
	assign a[WIDTH*150+:WIDTH]=-33670;
	assign a[WIDTH*151+:WIDTH]=50916;
	assign a[WIDTH*152+:WIDTH]=78914;
	assign a[WIDTH*153+:WIDTH]=29466;
	assign a[WIDTH*154+:WIDTH]=18865;
	assign a[WIDTH*155+:WIDTH]=43934;
	assign a[WIDTH*156+:WIDTH]=-50610;
	assign a[WIDTH*157+:WIDTH]=-7422;
	assign a[WIDTH*158+:WIDTH]=-64871;
	assign a[WIDTH*159+:WIDTH]=39927;
	assign a[WIDTH*160+:WIDTH]=42609;
	assign a[WIDTH*161+:WIDTH]=-2913;
	assign a[WIDTH*162+:WIDTH]=95817;
	assign a[WIDTH*163+:WIDTH]=-132556;
	assign a[WIDTH*164+:WIDTH]=-60073;
	assign a[WIDTH*165+:WIDTH]=-45502;
	assign a[WIDTH*166+:WIDTH]=87861;
	assign a[WIDTH*167+:WIDTH]=14700;
	assign a[WIDTH*168+:WIDTH]=41252;
	assign a[WIDTH*169+:WIDTH]=-77526;
	assign a[WIDTH*170+:WIDTH]=-91203;
	assign a[WIDTH*171+:WIDTH]=82734;
	assign a[WIDTH*172+:WIDTH]=77510;
	assign a[WIDTH*173+:WIDTH]=-99162;
	assign a[WIDTH*174+:WIDTH]=76605;
	assign a[WIDTH*175+:WIDTH]=51535;
	assign a[WIDTH*176+:WIDTH]=-145229;
	assign a[WIDTH*177+:WIDTH]=-23054;
	assign a[WIDTH*178+:WIDTH]=13348;
	assign a[WIDTH*179+:WIDTH]=75527;
	assign a[WIDTH*180+:WIDTH]=53485;
	assign a[WIDTH*181+:WIDTH]=-135533;
	assign a[WIDTH*182+:WIDTH]=-70671;
	assign a[WIDTH*183+:WIDTH]=85195;
	assign a[WIDTH*184+:WIDTH]=116404;
	assign a[WIDTH*185+:WIDTH]=164481;
	assign a[WIDTH*186+:WIDTH]=-41390;
	assign a[WIDTH*187+:WIDTH]=-61533;
	assign a[WIDTH*188+:WIDTH]=37731;
	assign a[WIDTH*189+:WIDTH]=79035;
	assign a[WIDTH*190+:WIDTH]=-31817;
	assign a[WIDTH*191+:WIDTH]=73314;
	assign a[WIDTH*192+:WIDTH]=-57535;
	assign a[WIDTH*193+:WIDTH]=141616;
	assign a[WIDTH*194+:WIDTH]=57235;
	assign a[WIDTH*195+:WIDTH]=-86884;
	assign a[WIDTH*196+:WIDTH]=-97992;
	assign a[WIDTH*197+:WIDTH]=67595;
	assign a[WIDTH*198+:WIDTH]=19962;
	assign a[WIDTH*199+:WIDTH]=-34643;
	assign a[WIDTH*200+:WIDTH]=15251;
	assign a[WIDTH*201+:WIDTH]=73229;
	assign a[WIDTH*202+:WIDTH]=-23620;
	assign a[WIDTH*203+:WIDTH]=45643;
	assign a[WIDTH*204+:WIDTH]=11508;
	assign a[WIDTH*205+:WIDTH]=3397;
	assign a[WIDTH*206+:WIDTH]=10189;
	assign a[WIDTH*207+:WIDTH]=-55406;
	assign a[WIDTH*208+:WIDTH]=13546;
	assign a[WIDTH*209+:WIDTH]=82506;
	assign a[WIDTH*210+:WIDTH]=81963;
	assign a[WIDTH*211+:WIDTH]=-71476;
	assign a[WIDTH*212+:WIDTH]=-22475;
	assign a[WIDTH*213+:WIDTH]=76258;
	assign a[WIDTH*214+:WIDTH]=-85306;
	assign a[WIDTH*215+:WIDTH]=-94963;
	assign a[WIDTH*216+:WIDTH]=-61251;
	assign a[WIDTH*217+:WIDTH]=21409;
	assign a[WIDTH*218+:WIDTH]=36340;
	assign a[WIDTH*219+:WIDTH]=42040;
	assign a[WIDTH*220+:WIDTH]=15541;
	assign a[WIDTH*221+:WIDTH]=114229;
	assign a[WIDTH*222+:WIDTH]=50381;
	assign a[WIDTH*223+:WIDTH]=-26741;
	assign a[WIDTH*224+:WIDTH]=25292;
	assign a[WIDTH*225+:WIDTH]=-24315;
	assign a[WIDTH*226+:WIDTH]=45830;
	assign a[WIDTH*227+:WIDTH]=71874;
	assign a[WIDTH*228+:WIDTH]=-89233;
	assign a[WIDTH*229+:WIDTH]=142732;
	assign a[WIDTH*230+:WIDTH]=47107;
	assign a[WIDTH*231+:WIDTH]=7566;
	assign a[WIDTH*232+:WIDTH]=22841;
	assign a[WIDTH*233+:WIDTH]=-179138;
	assign a[WIDTH*234+:WIDTH]=-56374;
	assign a[WIDTH*235+:WIDTH]=-8094;
	assign a[WIDTH*236+:WIDTH]=7890;
	assign a[WIDTH*237+:WIDTH]=52167;
	assign a[WIDTH*238+:WIDTH]=-85915;
	assign a[WIDTH*239+:WIDTH]=39728;
	assign a[WIDTH*240+:WIDTH]=10206;
	assign a[WIDTH*241+:WIDTH]=47191;
	assign a[WIDTH*242+:WIDTH]=50311;
	assign a[WIDTH*243+:WIDTH]=74375;
	assign a[WIDTH*244+:WIDTH]=-172028;
	assign a[WIDTH*245+:WIDTH]=17676;
	assign a[WIDTH*246+:WIDTH]=-45854;
	assign a[WIDTH*247+:WIDTH]=-63506;
	assign a[WIDTH*248+:WIDTH]=35449;
	assign a[WIDTH*249+:WIDTH]=-72229;
	assign a[WIDTH*250+:WIDTH]=6723;
	assign a[WIDTH*251+:WIDTH]=51821;
	assign a[WIDTH*252+:WIDTH]=-43760;
	assign a[WIDTH*253+:WIDTH]=-25921;
	assign a[WIDTH*254+:WIDTH]=22420;
	assign a[WIDTH*255+:WIDTH]=92223;
	assign a[WIDTH*256+:WIDTH]=-73775;
	assign a[WIDTH*257+:WIDTH]=-132268;
	assign a[WIDTH*258+:WIDTH]=115412;
	assign a[WIDTH*259+:WIDTH]=-58638;
	assign a[WIDTH*260+:WIDTH]=17003;
	assign a[WIDTH*261+:WIDTH]=9878;
	assign a[WIDTH*262+:WIDTH]=-49232;
	assign a[WIDTH*263+:WIDTH]=-34048;
	assign a[WIDTH*264+:WIDTH]=-7317;
	assign a[WIDTH*265+:WIDTH]=-83000;
	assign a[WIDTH*266+:WIDTH]=-104699;
	assign a[WIDTH*267+:WIDTH]=-7221;
	assign a[WIDTH*268+:WIDTH]=9695;
	assign a[WIDTH*269+:WIDTH]=19445;
	assign a[WIDTH*270+:WIDTH]=26904;
	assign a[WIDTH*271+:WIDTH]=70323;
	assign a[WIDTH*272+:WIDTH]=5358;
	assign a[WIDTH*273+:WIDTH]=75140;
	assign a[WIDTH*274+:WIDTH]=-68209;
	assign a[WIDTH*275+:WIDTH]=44693;
	assign a[WIDTH*276+:WIDTH]=-110049;
	assign a[WIDTH*277+:WIDTH]=-18915;
	assign a[WIDTH*278+:WIDTH]=80148;
	assign a[WIDTH*279+:WIDTH]=-11506;
	assign a[WIDTH*280+:WIDTH]=27558;
	assign a[WIDTH*281+:WIDTH]=9867;
	assign a[WIDTH*282+:WIDTH]=83727;
	assign a[WIDTH*283+:WIDTH]=61625;
	assign a[WIDTH*284+:WIDTH]=-65680;
	assign a[WIDTH*285+:WIDTH]=15675;
	assign a[WIDTH*286+:WIDTH]=66233;
	assign a[WIDTH*287+:WIDTH]=-100371;
	assign a[WIDTH*288+:WIDTH]=-59634;
	assign a[WIDTH*289+:WIDTH]=-18194;
	assign a[WIDTH*290+:WIDTH]=66391;
	assign a[WIDTH*291+:WIDTH]=-40501;
	assign a[WIDTH*292+:WIDTH]=9992;
	assign a[WIDTH*293+:WIDTH]=66078;
	assign a[WIDTH*294+:WIDTH]=-25654;
	assign a[WIDTH*295+:WIDTH]=30098;
	assign a[WIDTH*296+:WIDTH]=69724;
	assign a[WIDTH*297+:WIDTH]=65897;
	assign a[WIDTH*298+:WIDTH]=75042;
	assign a[WIDTH*299+:WIDTH]=-72830;
	assign a[WIDTH*300+:WIDTH]=8286;
	assign a[WIDTH*301+:WIDTH]=39488;
	assign a[WIDTH*302+:WIDTH]=106919;
	assign a[WIDTH*303+:WIDTH]=5375;
	assign a[WIDTH*304+:WIDTH]=106123;
	assign a[WIDTH*305+:WIDTH]=-81984;
	assign a[WIDTH*306+:WIDTH]=14189;
	assign a[WIDTH*307+:WIDTH]=80758;
	assign a[WIDTH*308+:WIDTH]=114153;
	assign a[WIDTH*309+:WIDTH]=49327;
	assign a[WIDTH*310+:WIDTH]=-78850;
	assign a[WIDTH*311+:WIDTH]=76112;
	assign a[WIDTH*312+:WIDTH]=-99904;
	assign a[WIDTH*313+:WIDTH]=-68179;
	assign a[WIDTH*314+:WIDTH]=42420;
	assign a[WIDTH*315+:WIDTH]=-143534;
	assign a[WIDTH*316+:WIDTH]=-64007;
	assign a[WIDTH*317+:WIDTH]=43160;
	assign a[WIDTH*318+:WIDTH]=104729;
	assign a[WIDTH*319+:WIDTH]=-58622;
	assign a[WIDTH*320+:WIDTH]=45040;
	assign a[WIDTH*321+:WIDTH]=104011;
	assign a[WIDTH*322+:WIDTH]=71271;
	assign a[WIDTH*323+:WIDTH]=59396;
	assign a[WIDTH*324+:WIDTH]=-101070;
	assign a[WIDTH*325+:WIDTH]=-20589;
	assign a[WIDTH*326+:WIDTH]=7275;
	assign a[WIDTH*327+:WIDTH]=73760;
	assign a[WIDTH*328+:WIDTH]=-15094;
	assign a[WIDTH*329+:WIDTH]=-18982;
	assign a[WIDTH*330+:WIDTH]=-71568;
	assign a[WIDTH*331+:WIDTH]=7772;
	assign a[WIDTH*332+:WIDTH]=-12390;
	assign a[WIDTH*333+:WIDTH]=8716;
	assign a[WIDTH*334+:WIDTH]=150140;
	assign a[WIDTH*335+:WIDTH]=25323;
	assign a[WIDTH*336+:WIDTH]=-6810;
	assign a[WIDTH*337+:WIDTH]=1295;
	assign a[WIDTH*338+:WIDTH]=134387;
	assign a[WIDTH*339+:WIDTH]=-52380;
	assign a[WIDTH*340+:WIDTH]=23535;
	assign a[WIDTH*341+:WIDTH]=-3096;
	assign a[WIDTH*342+:WIDTH]=-50652;
	assign a[WIDTH*343+:WIDTH]=84686;
	assign a[WIDTH*344+:WIDTH]=8683;
	assign a[WIDTH*345+:WIDTH]=13273;
	assign a[WIDTH*346+:WIDTH]=91716;
	assign a[WIDTH*347+:WIDTH]=-25270;
	assign a[WIDTH*348+:WIDTH]=-49575;
	assign a[WIDTH*349+:WIDTH]=-27001;
	assign a[WIDTH*350+:WIDTH]=-75782;
	assign a[WIDTH*351+:WIDTH]=26036;
	assign a[WIDTH*352+:WIDTH]=53432;
	assign a[WIDTH*353+:WIDTH]=-49904;
	assign a[WIDTH*354+:WIDTH]=-3338;
	assign a[WIDTH*355+:WIDTH]=14559;
	assign a[WIDTH*356+:WIDTH]=-18089;
	assign a[WIDTH*357+:WIDTH]=-80303;
	assign a[WIDTH*358+:WIDTH]=117004;
	assign a[WIDTH*359+:WIDTH]=108032;
	assign a[WIDTH*360+:WIDTH]=41109;
	assign a[WIDTH*361+:WIDTH]=-39178;
	assign a[WIDTH*362+:WIDTH]=-3384;
	assign a[WIDTH*363+:WIDTH]=-65671;
	assign a[WIDTH*364+:WIDTH]=68404;
	assign a[WIDTH*365+:WIDTH]=102236;
	assign a[WIDTH*366+:WIDTH]=-46783;
	assign a[WIDTH*367+:WIDTH]=-9150;
	assign a[WIDTH*368+:WIDTH]=6704;
	assign a[WIDTH*369+:WIDTH]=69992;
	assign a[WIDTH*370+:WIDTH]=74433;
	assign a[WIDTH*371+:WIDTH]=16568;
	assign a[WIDTH*372+:WIDTH]=-65220;
	assign a[WIDTH*373+:WIDTH]=-58860;
	assign a[WIDTH*374+:WIDTH]=-15762;
	assign a[WIDTH*375+:WIDTH]=-88042;
	assign a[WIDTH*376+:WIDTH]=-80821;
	assign a[WIDTH*377+:WIDTH]=-31866;
	assign a[WIDTH*378+:WIDTH]=-82747;
	assign a[WIDTH*379+:WIDTH]=-26198;
	assign a[WIDTH*380+:WIDTH]=-74575;
	assign a[WIDTH*381+:WIDTH]=30498;
	assign a[WIDTH*382+:WIDTH]=25076;
	assign a[WIDTH*383+:WIDTH]=-25411;
	assign a[WIDTH*384+:WIDTH]=-22372;
	assign a[WIDTH*385+:WIDTH]=64133;
	assign a[WIDTH*386+:WIDTH]=83206;
	assign a[WIDTH*387+:WIDTH]=60490;
	assign a[WIDTH*388+:WIDTH]=59171;
	assign a[WIDTH*389+:WIDTH]=35349;
	assign a[WIDTH*390+:WIDTH]=-5146;
	assign a[WIDTH*391+:WIDTH]=37739;
	assign a[WIDTH*392+:WIDTH]=-529;
	assign a[WIDTH*393+:WIDTH]=21373;
	assign a[WIDTH*394+:WIDTH]=25197;
	assign a[WIDTH*395+:WIDTH]=92272;
	assign a[WIDTH*396+:WIDTH]=-34018;
	assign a[WIDTH*397+:WIDTH]=47493;
	assign a[WIDTH*398+:WIDTH]=-93665;
	assign a[WIDTH*399+:WIDTH]=-38986;
	assign a[WIDTH*400+:WIDTH]=-46440;
	assign a[WIDTH*401+:WIDTH]=-41490;
	assign a[WIDTH*402+:WIDTH]=-3940;
	assign a[WIDTH*403+:WIDTH]=40057;
	assign a[WIDTH*404+:WIDTH]=115273;
	assign a[WIDTH*405+:WIDTH]=-108480;
	assign a[WIDTH*406+:WIDTH]=-91586;
	assign a[WIDTH*407+:WIDTH]=19014;
	assign a[WIDTH*408+:WIDTH]=-75089;
	assign a[WIDTH*409+:WIDTH]=31867;
	assign a[WIDTH*410+:WIDTH]=87194;
	assign a[WIDTH*411+:WIDTH]=63017;
	assign a[WIDTH*412+:WIDTH]=75833;
	assign a[WIDTH*413+:WIDTH]=70033;
	assign a[WIDTH*414+:WIDTH]=-77436;
	assign a[WIDTH*415+:WIDTH]=49899;
	assign a[WIDTH*416+:WIDTH]=-71157;
	assign a[WIDTH*417+:WIDTH]=51201;
	assign a[WIDTH*418+:WIDTH]=-77144;
	assign a[WIDTH*419+:WIDTH]=-6515;
	assign a[WIDTH*420+:WIDTH]=-30765;
	assign a[WIDTH*421+:WIDTH]=1480;
	assign a[WIDTH*422+:WIDTH]=161121;
	assign a[WIDTH*423+:WIDTH]=-148777;
	assign a[WIDTH*424+:WIDTH]=47802;
	assign a[WIDTH*425+:WIDTH]=182149;
	assign a[WIDTH*426+:WIDTH]=-33706;
	assign a[WIDTH*427+:WIDTH]=98043;
	assign a[WIDTH*428+:WIDTH]=49291;
	assign a[WIDTH*429+:WIDTH]=28391;
	assign a[WIDTH*430+:WIDTH]=69328;
	assign a[WIDTH*431+:WIDTH]=61419;
	assign a[WIDTH*432+:WIDTH]=-34649;
	assign a[WIDTH*433+:WIDTH]=-35910;
	assign a[WIDTH*434+:WIDTH]=36775;
	assign a[WIDTH*435+:WIDTH]=84485;
	assign a[WIDTH*436+:WIDTH]=14756;
	assign a[WIDTH*437+:WIDTH]=122566;
	assign a[WIDTH*438+:WIDTH]=-5500;
	assign a[WIDTH*439+:WIDTH]=79200;
	assign a[WIDTH*440+:WIDTH]=-72783;
	assign a[WIDTH*441+:WIDTH]=77974;
	assign a[WIDTH*442+:WIDTH]=67707;
	assign a[WIDTH*443+:WIDTH]=-62636;
	assign a[WIDTH*444+:WIDTH]=-75901;
	assign a[WIDTH*445+:WIDTH]=65800;
	assign a[WIDTH*446+:WIDTH]=-14979;
	assign a[WIDTH*447+:WIDTH]=-54276;
	assign a[WIDTH*448+:WIDTH]=52262;
	assign a[WIDTH*449+:WIDTH]=3940;
	assign a[WIDTH*450+:WIDTH]=14138;
	assign a[WIDTH*451+:WIDTH]=16012;
	assign a[WIDTH*452+:WIDTH]=-29179;
	assign a[WIDTH*453+:WIDTH]=56617;
	assign a[WIDTH*454+:WIDTH]=-53911;
	assign a[WIDTH*455+:WIDTH]=-45151;
	assign a[WIDTH*456+:WIDTH]=51013;
	assign a[WIDTH*457+:WIDTH]=76349;
	assign a[WIDTH*458+:WIDTH]=35985;
	assign a[WIDTH*459+:WIDTH]=89348;
	assign a[WIDTH*460+:WIDTH]=-26399;
	assign a[WIDTH*461+:WIDTH]=-62111;
	assign a[WIDTH*462+:WIDTH]=26295;
	assign a[WIDTH*463+:WIDTH]=147447;
	assign a[WIDTH*464+:WIDTH]=-123761;
	assign a[WIDTH*465+:WIDTH]=-118817;
	assign a[WIDTH*466+:WIDTH]=-99903;
	assign a[WIDTH*467+:WIDTH]=-55444;
	assign a[WIDTH*468+:WIDTH]=79075;
	assign a[WIDTH*469+:WIDTH]=24275;
	assign a[WIDTH*470+:WIDTH]=-158533;
	assign a[WIDTH*471+:WIDTH]=-22772;
	assign a[WIDTH*472+:WIDTH]=-41062;
	assign a[WIDTH*473+:WIDTH]=29262;
	assign a[WIDTH*474+:WIDTH]=-121788;
	assign a[WIDTH*475+:WIDTH]=-93031;
	assign a[WIDTH*476+:WIDTH]=4123;
	assign a[WIDTH*477+:WIDTH]=5167;
	assign a[WIDTH*478+:WIDTH]=-8994;
	assign a[WIDTH*479+:WIDTH]=7067;
	assign a[WIDTH*480+:WIDTH]=37358;
	assign a[WIDTH*481+:WIDTH]=-48873;
	assign a[WIDTH*482+:WIDTH]=11033;
	assign a[WIDTH*483+:WIDTH]=-68925;
	assign a[WIDTH*484+:WIDTH]=7168;
	assign a[WIDTH*485+:WIDTH]=37270;
	assign a[WIDTH*486+:WIDTH]=-53423;
	assign a[WIDTH*487+:WIDTH]=-38850;
	assign a[WIDTH*488+:WIDTH]=-26521;
	assign a[WIDTH*489+:WIDTH]=89514;
	assign a[WIDTH*490+:WIDTH]=-7784;
	assign a[WIDTH*491+:WIDTH]=3394;
	assign a[WIDTH*492+:WIDTH]=-26210;
	assign a[WIDTH*493+:WIDTH]=-2230;
	assign a[WIDTH*494+:WIDTH]=-74265;
	assign a[WIDTH*495+:WIDTH]=66176;
	assign a[WIDTH*496+:WIDTH]=-152457;
	assign a[WIDTH*497+:WIDTH]=12254;
	assign a[WIDTH*498+:WIDTH]=4701;
	assign a[WIDTH*499+:WIDTH]=-110129;
	assign a[WIDTH*500+:WIDTH]=14186;
	assign a[WIDTH*501+:WIDTH]=21983;
	assign a[WIDTH*502+:WIDTH]=57939;
	assign a[WIDTH*503+:WIDTH]=-55634;
	assign a[WIDTH*504+:WIDTH]=-36282;
	assign a[WIDTH*505+:WIDTH]=-89092;
	assign a[WIDTH*506+:WIDTH]=68086;
	assign a[WIDTH*507+:WIDTH]=-44312;
	assign a[WIDTH*508+:WIDTH]=11293;
	assign a[WIDTH*509+:WIDTH]=-6124;
	assign a[WIDTH*510+:WIDTH]=-70185;
	assign a[WIDTH*511+:WIDTH]=112626;

endmodule
