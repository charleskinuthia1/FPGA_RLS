`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   12:42:35 03/31/2016
// Design Name:   RLS
// Module Name:   C:/Users/Charlz/Documents/3_KTH/KEX_Xillinc/RLS/RLS_tb.v
// Project Name:  RLS
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: RLS
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module RLS_tb;
	parameter WIDTH=32;
	parameter SIZE=16;
	parameter ITER=32;
	parameter COMBSIZE = 4;
	
	// Inputs
	reg clk;
	reg reset;
	reg [SIZE*WIDTH-1:0] x0;
	reg [SIZE*ITER*WIDTH-1:0] k;
	reg [ITER*WIDTH-1:0] b;
	reg [SIZE*ITER*WIDTH-1:0] a;

	// Outputs
	wire [SIZE*WIDTH-1:0] x;
	wire ready;

	// Instantiate the Unit Under Test (UUT)
	RLSBlock #(.WIDTH(WIDTH), .SIZE(SIZE),.ITER(ITER), .COMBSIZE(COMBSIZE)) uut (
		.clk(clk), 
		.reset(reset), 
		.x0(x0), 
		.k_SIZE(k), 
		.b_SIZE(b), 
		.a_SIZE(a), 
		.x(x), 
		.ready(ready)
	);
	
	always begin
		#15 clk=~clk;
	end
	
	task nextData;
	begin
		k <= k>>WIDTH*ITER;
	end
	endtask;
	
	task initk;
	begin
	k[WIDTH*0+:WIDTH]=2.0**16*-0.00675739;
k[WIDTH*1+:WIDTH]=2.0**16*-0.11864723;
k[WIDTH*2+:WIDTH]=2.0**16*0.10293554;
k[WIDTH*3+:WIDTH]=2.0**16*0.01747938;
k[WIDTH*4+:WIDTH]=2.0**16*0.03989958;
k[WIDTH*5+:WIDTH]=2.0**16*-0.00380982;
k[WIDTH*6+:WIDTH]=2.0**16*-0.01201210;
k[WIDTH*7+:WIDTH]=2.0**16*-0.11122228;
k[WIDTH*8+:WIDTH]=2.0**16*0.11480459;
k[WIDTH*9+:WIDTH]=2.0**16*0.07711716;
k[WIDTH*10+:WIDTH]=2.0**16*-0.07760189;
k[WIDTH*11+:WIDTH]=2.0**16*-0.01708212;
k[WIDTH*12+:WIDTH]=2.0**16*-0.07820042;
k[WIDTH*13+:WIDTH]=2.0**16*-0.03163632;
k[WIDTH*14+:WIDTH]=2.0**16*-0.00728598;
k[WIDTH*15+:WIDTH]=2.0**16*0.04311193;
k[WIDTH*16+:WIDTH]=2.0**16*0.12380668;
k[WIDTH*17+:WIDTH]=2.0**16*-0.01953538;
k[WIDTH*18+:WIDTH]=2.0**16*-0.00241381;
k[WIDTH*19+:WIDTH]=2.0**16*-0.04492235;
k[WIDTH*20+:WIDTH]=2.0**16*-0.05669642;
k[WIDTH*21+:WIDTH]=2.0**16*-0.03005831;
k[WIDTH*22+:WIDTH]=2.0**16*-0.00345552;
k[WIDTH*23+:WIDTH]=2.0**16*-0.02821819;
k[WIDTH*24+:WIDTH]=2.0**16*-0.06521373;
k[WIDTH*25+:WIDTH]=2.0**16*-0.06318049;
k[WIDTH*26+:WIDTH]=2.0**16*-0.05835912;
k[WIDTH*27+:WIDTH]=2.0**16*-0.08560921;
k[WIDTH*28+:WIDTH]=2.0**16*0.02709743;
k[WIDTH*29+:WIDTH]=2.0**16*-0.04897373;
k[WIDTH*30+:WIDTH]=2.0**16*0.01725284;
k[WIDTH*31+:WIDTH]=2.0**16*0.00982406;
k[WIDTH*32+:WIDTH]=2.0**16*-0.10797052;
k[WIDTH*33+:WIDTH]=2.0**16*-0.10678354;
k[WIDTH*34+:WIDTH]=2.0**16*-0.06378132;
k[WIDTH*35+:WIDTH]=2.0**16*-0.02485593;
k[WIDTH*36+:WIDTH]=2.0**16*-0.02192487;
k[WIDTH*37+:WIDTH]=2.0**16*-0.05023058;
k[WIDTH*38+:WIDTH]=2.0**16*-0.00435302;
k[WIDTH*39+:WIDTH]=2.0**16*-0.02312640;
k[WIDTH*40+:WIDTH]=2.0**16*0.05547411;
k[WIDTH*41+:WIDTH]=2.0**16*-0.03333542;
k[WIDTH*42+:WIDTH]=2.0**16*-0.02953023;
k[WIDTH*43+:WIDTH]=2.0**16*0.04860764;
k[WIDTH*44+:WIDTH]=2.0**16*0.05629476;
k[WIDTH*45+:WIDTH]=2.0**16*-0.00898510;
k[WIDTH*46+:WIDTH]=2.0**16*0.00497664;
k[WIDTH*47+:WIDTH]=2.0**16*-0.00899659;
k[WIDTH*48+:WIDTH]=2.0**16*0.01284226;
k[WIDTH*49+:WIDTH]=2.0**16*0.04990850;
k[WIDTH*50+:WIDTH]=2.0**16*-0.02493618;
k[WIDTH*51+:WIDTH]=2.0**16*-0.08680240;
k[WIDTH*52+:WIDTH]=2.0**16*-0.04665895;
k[WIDTH*53+:WIDTH]=2.0**16*0.12318097;
k[WIDTH*54+:WIDTH]=2.0**16*0.02577212;
k[WIDTH*55+:WIDTH]=2.0**16*-0.00682386;
k[WIDTH*56+:WIDTH]=2.0**16*0.08354079;
k[WIDTH*57+:WIDTH]=2.0**16*-0.05108302;
k[WIDTH*58+:WIDTH]=2.0**16*0.00464850;
k[WIDTH*59+:WIDTH]=2.0**16*0.00630319;
k[WIDTH*60+:WIDTH]=2.0**16*0.01060614;
k[WIDTH*61+:WIDTH]=2.0**16*-0.04071465;
k[WIDTH*62+:WIDTH]=2.0**16*-0.08004992;
k[WIDTH*63+:WIDTH]=2.0**16*0.05954602;
k[WIDTH*64+:WIDTH]=2.0**16*0.09988593;
k[WIDTH*65+:WIDTH]=2.0**16*-0.04225802;
k[WIDTH*66+:WIDTH]=2.0**16*-0.14288966;
k[WIDTH*67+:WIDTH]=2.0**16*0.18961658;
k[WIDTH*68+:WIDTH]=2.0**16*-0.17202424;
k[WIDTH*69+:WIDTH]=2.0**16*0.00874481;
k[WIDTH*70+:WIDTH]=2.0**16*0.05207024;
k[WIDTH*71+:WIDTH]=2.0**16*-0.01726722;
k[WIDTH*72+:WIDTH]=2.0**16*0.00598238;
k[WIDTH*73+:WIDTH]=2.0**16*0.09388509;
k[WIDTH*74+:WIDTH]=2.0**16*-0.00383367;
k[WIDTH*75+:WIDTH]=2.0**16*-0.03546520;
k[WIDTH*76+:WIDTH]=2.0**16*-0.04286238;
k[WIDTH*77+:WIDTH]=2.0**16*-0.06535106;
k[WIDTH*78+:WIDTH]=2.0**16*-0.03690350;
k[WIDTH*79+:WIDTH]=2.0**16*0.09092682;
k[WIDTH*80+:WIDTH]=2.0**16*-0.10788038;
k[WIDTH*81+:WIDTH]=2.0**16*-0.03878917;
k[WIDTH*82+:WIDTH]=2.0**16*0.14796845;
k[WIDTH*83+:WIDTH]=2.0**16*-0.12177139;
k[WIDTH*84+:WIDTH]=2.0**16*-0.01770701;
k[WIDTH*85+:WIDTH]=2.0**16*0.10670917;
k[WIDTH*86+:WIDTH]=2.0**16*0.03036475;
k[WIDTH*87+:WIDTH]=2.0**16*0.01113235;
k[WIDTH*88+:WIDTH]=2.0**16*-0.08303959;
k[WIDTH*89+:WIDTH]=2.0**16*0.12595029;
k[WIDTH*90+:WIDTH]=2.0**16*0.09038787;
k[WIDTH*91+:WIDTH]=2.0**16*0.03061880;
k[WIDTH*92+:WIDTH]=2.0**16*0.02590304;
k[WIDTH*93+:WIDTH]=2.0**16*-0.05492817;
k[WIDTH*94+:WIDTH]=2.0**16*0.01440852;
k[WIDTH*95+:WIDTH]=2.0**16*-0.00865741;
k[WIDTH*96+:WIDTH]=2.0**16*-0.19220649;
k[WIDTH*97+:WIDTH]=2.0**16*0.09177092;
k[WIDTH*98+:WIDTH]=2.0**16*-0.10008910;
k[WIDTH*99+:WIDTH]=2.0**16*-0.11025599;
k[WIDTH*100+:WIDTH]=2.0**16*-0.01771940;
k[WIDTH*101+:WIDTH]=2.0**16*-0.16833076;
k[WIDTH*102+:WIDTH]=2.0**16*0.04380171;
k[WIDTH*103+:WIDTH]=2.0**16*0.08003279;
k[WIDTH*104+:WIDTH]=2.0**16*-0.10295565;
k[WIDTH*105+:WIDTH]=2.0**16*0.02511828;
k[WIDTH*106+:WIDTH]=2.0**16*-0.31061323;
k[WIDTH*107+:WIDTH]=2.0**16*-0.05572486;
k[WIDTH*108+:WIDTH]=2.0**16*-0.19247220;
k[WIDTH*109+:WIDTH]=2.0**16*-0.10028265;
k[WIDTH*110+:WIDTH]=2.0**16*-0.00810042;
k[WIDTH*111+:WIDTH]=2.0**16*0.16322996;
k[WIDTH*112+:WIDTH]=2.0**16*0.02568036;
k[WIDTH*113+:WIDTH]=2.0**16*-0.08255348;
k[WIDTH*114+:WIDTH]=2.0**16*0.03726446;
k[WIDTH*115+:WIDTH]=2.0**16*0.05428324;
k[WIDTH*116+:WIDTH]=2.0**16*0.05822590;
k[WIDTH*117+:WIDTH]=2.0**16*-0.13969586;
k[WIDTH*118+:WIDTH]=2.0**16*0.27549265;
k[WIDTH*119+:WIDTH]=2.0**16*-0.13654676;
k[WIDTH*120+:WIDTH]=2.0**16*-0.11249848;
k[WIDTH*121+:WIDTH]=2.0**16*-0.17639137;
k[WIDTH*122+:WIDTH]=2.0**16*0.06430571;
k[WIDTH*123+:WIDTH]=2.0**16*0.05855291;
k[WIDTH*124+:WIDTH]=2.0**16*-0.14681439;
k[WIDTH*125+:WIDTH]=2.0**16*0.16080800;
k[WIDTH*126+:WIDTH]=2.0**16*-0.28455197;
k[WIDTH*127+:WIDTH]=2.0**16*-0.17371690;
k[WIDTH*128+:WIDTH]=2.0**16*0.08280505;
k[WIDTH*129+:WIDTH]=2.0**16*-0.05178405;
k[WIDTH*130+:WIDTH]=2.0**16*0.07377107;
k[WIDTH*131+:WIDTH]=2.0**16*0.03954268;
k[WIDTH*132+:WIDTH]=2.0**16*-0.03964575;
k[WIDTH*133+:WIDTH]=2.0**16*0.02120091;
k[WIDTH*134+:WIDTH]=2.0**16*0.06107968;
k[WIDTH*135+:WIDTH]=2.0**16*-0.00288359;
k[WIDTH*136+:WIDTH]=2.0**16*-0.00877551;
k[WIDTH*137+:WIDTH]=2.0**16*-0.16993842;
k[WIDTH*138+:WIDTH]=2.0**16*-0.11102028;
k[WIDTH*139+:WIDTH]=2.0**16*0.17713787;
k[WIDTH*140+:WIDTH]=2.0**16*-0.11760237;
k[WIDTH*141+:WIDTH]=2.0**16*0.04656787;
k[WIDTH*142+:WIDTH]=2.0**16*0.06398774;
k[WIDTH*143+:WIDTH]=2.0**16*0.02203650;
k[WIDTH*144+:WIDTH]=2.0**16*0.12542026;
k[WIDTH*145+:WIDTH]=2.0**16*-0.06505370;
k[WIDTH*146+:WIDTH]=2.0**16*-0.06987229;
k[WIDTH*147+:WIDTH]=2.0**16*-0.15973105;
k[WIDTH*148+:WIDTH]=2.0**16*0.03717368;
k[WIDTH*149+:WIDTH]=2.0**16*0.00416851;
k[WIDTH*150+:WIDTH]=2.0**16*-0.14173909;
k[WIDTH*151+:WIDTH]=2.0**16*0.01809618;
k[WIDTH*152+:WIDTH]=2.0**16*-0.06171712;
k[WIDTH*153+:WIDTH]=2.0**16*0.06660571;
k[WIDTH*154+:WIDTH]=2.0**16*0.09926338;
k[WIDTH*155+:WIDTH]=2.0**16*0.10735105;
k[WIDTH*156+:WIDTH]=2.0**16*-0.11423135;
k[WIDTH*157+:WIDTH]=2.0**16*0.02164126;
k[WIDTH*158+:WIDTH]=2.0**16*-0.02432526;
k[WIDTH*159+:WIDTH]=2.0**16*0.14632648;
k[WIDTH*160+:WIDTH]=2.0**16*-0.07174021;
k[WIDTH*161+:WIDTH]=2.0**16*0.20552124;
k[WIDTH*162+:WIDTH]=2.0**16*0.02790155;
k[WIDTH*163+:WIDTH]=2.0**16*-0.18916687;
k[WIDTH*164+:WIDTH]=2.0**16*-0.06256805;
k[WIDTH*165+:WIDTH]=2.0**16*-0.03377220;
k[WIDTH*166+:WIDTH]=2.0**16*0.09552039;
k[WIDTH*167+:WIDTH]=2.0**16*-0.35913331;
k[WIDTH*168+:WIDTH]=2.0**16*0.05615996;
k[WIDTH*169+:WIDTH]=2.0**16*-0.01216300;
k[WIDTH*170+:WIDTH]=2.0**16*0.11826205;
k[WIDTH*171+:WIDTH]=2.0**16*0.10862434;
k[WIDTH*172+:WIDTH]=2.0**16*0.06651045;
k[WIDTH*173+:WIDTH]=2.0**16*0.36067600;
k[WIDTH*174+:WIDTH]=2.0**16*0.06316681;
k[WIDTH*175+:WIDTH]=2.0**16*0.05587686;
k[WIDTH*176+:WIDTH]=2.0**16*-0.01095386;
k[WIDTH*177+:WIDTH]=2.0**16*-0.04073698;
k[WIDTH*178+:WIDTH]=2.0**16*-0.08701058;
k[WIDTH*179+:WIDTH]=2.0**16*0.09418784;
k[WIDTH*180+:WIDTH]=2.0**16*0.30264858;
k[WIDTH*181+:WIDTH]=2.0**16*0.01093193;
k[WIDTH*182+:WIDTH]=2.0**16*0.30870163;
k[WIDTH*183+:WIDTH]=2.0**16*-0.11929776;
k[WIDTH*184+:WIDTH]=2.0**16*-0.00746429;
k[WIDTH*185+:WIDTH]=2.0**16*-0.18582569;
k[WIDTH*186+:WIDTH]=2.0**16*-0.01096193;
k[WIDTH*187+:WIDTH]=2.0**16*-0.09125229;
k[WIDTH*188+:WIDTH]=2.0**16*0.01459386;
k[WIDTH*189+:WIDTH]=2.0**16*-0.21540690;
k[WIDTH*190+:WIDTH]=2.0**16*0.30872840;
k[WIDTH*191+:WIDTH]=2.0**16*0.20770746;
k[WIDTH*192+:WIDTH]=2.0**16*0.05436220;
k[WIDTH*193+:WIDTH]=2.0**16*-0.12879999;
k[WIDTH*194+:WIDTH]=2.0**16*-0.02088379;
k[WIDTH*195+:WIDTH]=2.0**16*-0.14230399;
k[WIDTH*196+:WIDTH]=2.0**16*0.05191997;
k[WIDTH*197+:WIDTH]=2.0**16*-0.04316867;
k[WIDTH*198+:WIDTH]=2.0**16*0.04496560;
k[WIDTH*199+:WIDTH]=2.0**16*0.35177427;
k[WIDTH*200+:WIDTH]=2.0**16*0.06717479;
k[WIDTH*201+:WIDTH]=2.0**16*0.12062075;
k[WIDTH*202+:WIDTH]=2.0**16*-0.01330731;
k[WIDTH*203+:WIDTH]=2.0**16*-0.18694566;
k[WIDTH*204+:WIDTH]=2.0**16*0.09401296;
k[WIDTH*205+:WIDTH]=2.0**16*0.51316289;
k[WIDTH*206+:WIDTH]=2.0**16*-0.10775499;
k[WIDTH*207+:WIDTH]=2.0**16*0.36070573;
k[WIDTH*208+:WIDTH]=2.0**16*-0.09639928;
k[WIDTH*209+:WIDTH]=2.0**16*-0.01970282;
k[WIDTH*210+:WIDTH]=2.0**16*-0.06919518;
k[WIDTH*211+:WIDTH]=2.0**16*0.09357052;
k[WIDTH*212+:WIDTH]=2.0**16*0.09692758;
k[WIDTH*213+:WIDTH]=2.0**16*0.13048034;
k[WIDTH*214+:WIDTH]=2.0**16*-0.02609143;
k[WIDTH*215+:WIDTH]=2.0**16*-0.24361973;
k[WIDTH*216+:WIDTH]=2.0**16*-0.10282420;
k[WIDTH*217+:WIDTH]=2.0**16*-0.00547956;
k[WIDTH*218+:WIDTH]=2.0**16*-0.13174015;
k[WIDTH*219+:WIDTH]=2.0**16*-0.01731902;
k[WIDTH*220+:WIDTH]=2.0**16*0.15246645;
k[WIDTH*221+:WIDTH]=2.0**16*0.07286580;
k[WIDTH*222+:WIDTH]=2.0**16*0.05933490;
k[WIDTH*223+:WIDTH]=2.0**16*0.18749520;
k[WIDTH*224+:WIDTH]=2.0**16*0.02603851;
k[WIDTH*225+:WIDTH]=2.0**16*0.09996840;
k[WIDTH*226+:WIDTH]=2.0**16*0.09871121;
k[WIDTH*227+:WIDTH]=2.0**16*-0.12265299;
k[WIDTH*228+:WIDTH]=2.0**16*-0.03559634;
k[WIDTH*229+:WIDTH]=2.0**16*-0.11531837;
k[WIDTH*230+:WIDTH]=2.0**16*0.04568064;
k[WIDTH*231+:WIDTH]=2.0**16*-0.02153681;
k[WIDTH*232+:WIDTH]=2.0**16*0.12374873;
k[WIDTH*233+:WIDTH]=2.0**16*0.02432216;
k[WIDTH*234+:WIDTH]=2.0**16*0.12778560;
k[WIDTH*235+:WIDTH]=2.0**16*-0.00536436;
k[WIDTH*236+:WIDTH]=2.0**16*0.14135647;
k[WIDTH*237+:WIDTH]=2.0**16*0.22507661;
k[WIDTH*238+:WIDTH]=2.0**16*0.02591619;
k[WIDTH*239+:WIDTH]=2.0**16*0.31092909;
k[WIDTH*240+:WIDTH]=2.0**16*0.04440602;
k[WIDTH*241+:WIDTH]=2.0**16*-0.07463081;
k[WIDTH*242+:WIDTH]=2.0**16*-0.27988326;
k[WIDTH*243+:WIDTH]=2.0**16*-0.32739451;
k[WIDTH*244+:WIDTH]=2.0**16*0.11501872;
k[WIDTH*245+:WIDTH]=2.0**16*0.19402599;
k[WIDTH*246+:WIDTH]=2.0**16*0.18881082;
k[WIDTH*247+:WIDTH]=2.0**16*0.13615659;
k[WIDTH*248+:WIDTH]=2.0**16*0.02956528;
k[WIDTH*249+:WIDTH]=2.0**16*0.19373246;
k[WIDTH*250+:WIDTH]=2.0**16*-0.26592240;
k[WIDTH*251+:WIDTH]=2.0**16*-0.12616829;
k[WIDTH*252+:WIDTH]=2.0**16*-0.18837504;
k[WIDTH*253+:WIDTH]=2.0**16*0.21153999;
k[WIDTH*254+:WIDTH]=2.0**16*0.23878130;
k[WIDTH*255+:WIDTH]=2.0**16*-0.38150082;
k[WIDTH*256+:WIDTH]=2.0**16*0.06814217;
k[WIDTH*257+:WIDTH]=2.0**16*0.10773576;
k[WIDTH*258+:WIDTH]=2.0**16*0.08531464;
k[WIDTH*259+:WIDTH]=2.0**16*0.05513094;
k[WIDTH*260+:WIDTH]=2.0**16*-0.06563171;
k[WIDTH*261+:WIDTH]=2.0**16*-0.10965987;
k[WIDTH*262+:WIDTH]=2.0**16*-0.01630461;
k[WIDTH*263+:WIDTH]=2.0**16*-0.06339886;
k[WIDTH*264+:WIDTH]=2.0**16*0.05091481;
k[WIDTH*265+:WIDTH]=2.0**16*0.04090749;
k[WIDTH*266+:WIDTH]=2.0**16*0.10897283;
k[WIDTH*267+:WIDTH]=2.0**16*0.08715862;
k[WIDTH*268+:WIDTH]=2.0**16*0.13493898;
k[WIDTH*269+:WIDTH]=2.0**16*-0.00748847;
k[WIDTH*270+:WIDTH]=2.0**16*-0.09784443;
k[WIDTH*271+:WIDTH]=2.0**16*-0.04161748;
k[WIDTH*272+:WIDTH]=2.0**16*0.12803741;
k[WIDTH*273+:WIDTH]=2.0**16*0.07573995;
k[WIDTH*274+:WIDTH]=2.0**16*-0.04143147;
k[WIDTH*275+:WIDTH]=2.0**16*-0.17295507;
k[WIDTH*276+:WIDTH]=2.0**16*-0.05792705;
k[WIDTH*277+:WIDTH]=2.0**16*-0.05684038;
k[WIDTH*278+:WIDTH]=2.0**16*0.14012211;
k[WIDTH*279+:WIDTH]=2.0**16*0.02179145;
k[WIDTH*280+:WIDTH]=2.0**16*0.04231609;
k[WIDTH*281+:WIDTH]=2.0**16*0.10981104;
k[WIDTH*282+:WIDTH]=2.0**16*0.03160763;
k[WIDTH*283+:WIDTH]=2.0**16*0.14867193;
k[WIDTH*284+:WIDTH]=2.0**16*-0.11023922;
k[WIDTH*285+:WIDTH]=2.0**16*-0.04187044;
k[WIDTH*286+:WIDTH]=2.0**16*0.04476972;
k[WIDTH*287+:WIDTH]=2.0**16*-0.32021851;
k[WIDTH*288+:WIDTH]=2.0**16*-0.08086230;
k[WIDTH*289+:WIDTH]=2.0**16*-0.02065023;
k[WIDTH*290+:WIDTH]=2.0**16*0.05444043;
k[WIDTH*291+:WIDTH]=2.0**16*0.02183418;
k[WIDTH*292+:WIDTH]=2.0**16*-0.17219796;
k[WIDTH*293+:WIDTH]=2.0**16*-0.02336010;
k[WIDTH*294+:WIDTH]=2.0**16*-0.17408705;
k[WIDTH*295+:WIDTH]=2.0**16*0.02851014;
k[WIDTH*296+:WIDTH]=2.0**16*-0.02954879;
k[WIDTH*297+:WIDTH]=2.0**16*-0.11048806;
k[WIDTH*298+:WIDTH]=2.0**16*0.02533973;
k[WIDTH*299+:WIDTH]=2.0**16*0.01703139;
k[WIDTH*300+:WIDTH]=2.0**16*-0.25169327;
k[WIDTH*301+:WIDTH]=2.0**16*-0.21289275;
k[WIDTH*302+:WIDTH]=2.0**16*-0.00041118;
k[WIDTH*303+:WIDTH]=2.0**16*-0.02084689;
k[WIDTH*304+:WIDTH]=2.0**16*0.02148715;
k[WIDTH*305+:WIDTH]=2.0**16*0.01343004;
k[WIDTH*306+:WIDTH]=2.0**16*0.11922884;
k[WIDTH*307+:WIDTH]=2.0**16*-0.05824952;
k[WIDTH*308+:WIDTH]=2.0**16*-0.03781781;
k[WIDTH*309+:WIDTH]=2.0**16*-0.08071795;
k[WIDTH*310+:WIDTH]=2.0**16*0.14365429;
k[WIDTH*311+:WIDTH]=2.0**16*0.11706908;
k[WIDTH*312+:WIDTH]=2.0**16*0.12103990;
k[WIDTH*313+:WIDTH]=2.0**16*-0.12443966;
k[WIDTH*314+:WIDTH]=2.0**16*0.16756184;
k[WIDTH*315+:WIDTH]=2.0**16*-0.00430685;
k[WIDTH*316+:WIDTH]=2.0**16*-0.17012493;
k[WIDTH*317+:WIDTH]=2.0**16*-0.10945135;
k[WIDTH*318+:WIDTH]=2.0**16*0.14905171;
k[WIDTH*319+:WIDTH]=2.0**16*0.07104986;
k[WIDTH*320+:WIDTH]=2.0**16*-0.04622265;
k[WIDTH*321+:WIDTH]=2.0**16*-0.01424641;
k[WIDTH*322+:WIDTH]=2.0**16*-0.06234612;
k[WIDTH*323+:WIDTH]=2.0**16*0.02495415;
k[WIDTH*324+:WIDTH]=2.0**16*-0.13200357;
k[WIDTH*325+:WIDTH]=2.0**16*0.03414088;
k[WIDTH*326+:WIDTH]=2.0**16*-0.10623316;
k[WIDTH*327+:WIDTH]=2.0**16*-0.06569616;
k[WIDTH*328+:WIDTH]=2.0**16*-0.10226254;
k[WIDTH*329+:WIDTH]=2.0**16*0.03520991;
k[WIDTH*330+:WIDTH]=2.0**16*-0.02975866;
k[WIDTH*331+:WIDTH]=2.0**16*0.04148075;
k[WIDTH*332+:WIDTH]=2.0**16*-0.09040951;
k[WIDTH*333+:WIDTH]=2.0**16*-0.05611680;
k[WIDTH*334+:WIDTH]=2.0**16*0.00043692;
k[WIDTH*335+:WIDTH]=2.0**16*-0.11068864;
k[WIDTH*336+:WIDTH]=2.0**16*-0.11740855;
k[WIDTH*337+:WIDTH]=2.0**16*-0.03695129;
k[WIDTH*338+:WIDTH]=2.0**16*0.00764025;
k[WIDTH*339+:WIDTH]=2.0**16*-0.08493642;
k[WIDTH*340+:WIDTH]=2.0**16*-0.04661258;
k[WIDTH*341+:WIDTH]=2.0**16*0.03831233;
k[WIDTH*342+:WIDTH]=2.0**16*-0.10744305;
k[WIDTH*343+:WIDTH]=2.0**16*-0.03555984;
k[WIDTH*344+:WIDTH]=2.0**16*0.03929477;
k[WIDTH*345+:WIDTH]=2.0**16*-0.12752402;
k[WIDTH*346+:WIDTH]=2.0**16*0.09866019;
k[WIDTH*347+:WIDTH]=2.0**16*-0.14635170;
k[WIDTH*348+:WIDTH]=2.0**16*-0.19330478;
k[WIDTH*349+:WIDTH]=2.0**16*0.04706220;
k[WIDTH*350+:WIDTH]=2.0**16*0.10830507;
k[WIDTH*351+:WIDTH]=2.0**16*0.07241234;
k[WIDTH*352+:WIDTH]=2.0**16*0.11430179;
k[WIDTH*353+:WIDTH]=2.0**16*0.02778084;
k[WIDTH*354+:WIDTH]=2.0**16*0.02904756;
k[WIDTH*355+:WIDTH]=2.0**16*0.05734162;
k[WIDTH*356+:WIDTH]=2.0**16*0.07841838;
k[WIDTH*357+:WIDTH]=2.0**16*-0.03876360;
k[WIDTH*358+:WIDTH]=2.0**16*0.04921332;
k[WIDTH*359+:WIDTH]=2.0**16*-0.00606343;
k[WIDTH*360+:WIDTH]=2.0**16*-0.04528686;
k[WIDTH*361+:WIDTH]=2.0**16*0.17084286;
k[WIDTH*362+:WIDTH]=2.0**16*-0.15827069;
k[WIDTH*363+:WIDTH]=2.0**16*0.15009844;
k[WIDTH*364+:WIDTH]=2.0**16*0.28879574;
k[WIDTH*365+:WIDTH]=2.0**16*0.04899369;
k[WIDTH*366+:WIDTH]=2.0**16*-0.13397305;
k[WIDTH*367+:WIDTH]=2.0**16*0.05235837;
k[WIDTH*368+:WIDTH]=2.0**16*-0.00039815;
k[WIDTH*369+:WIDTH]=2.0**16*0.04490141;
k[WIDTH*370+:WIDTH]=2.0**16*0.04415771;
k[WIDTH*371+:WIDTH]=2.0**16*-0.06910418;
k[WIDTH*372+:WIDTH]=2.0**16*-0.04277270;
k[WIDTH*373+:WIDTH]=2.0**16*-0.08593121;
k[WIDTH*374+:WIDTH]=2.0**16*-0.06989283;
k[WIDTH*375+:WIDTH]=2.0**16*0.07209670;
k[WIDTH*376+:WIDTH]=2.0**16*0.10410604;
k[WIDTH*377+:WIDTH]=2.0**16*-0.08987896;
k[WIDTH*378+:WIDTH]=2.0**16*0.12607388;
k[WIDTH*379+:WIDTH]=2.0**16*-0.02756430;
k[WIDTH*380+:WIDTH]=2.0**16*-0.10688521;
k[WIDTH*381+:WIDTH]=2.0**16*-0.04219642;
k[WIDTH*382+:WIDTH]=2.0**16*0.10363740;
k[WIDTH*383+:WIDTH]=2.0**16*0.08166745;
k[WIDTH*384+:WIDTH]=2.0**16*-0.01538773;
k[WIDTH*385+:WIDTH]=2.0**16*-0.06911971;
k[WIDTH*386+:WIDTH]=2.0**16*0.06497358;
k[WIDTH*387+:WIDTH]=2.0**16*0.11981118;
k[WIDTH*388+:WIDTH]=2.0**16*-0.01376406;
k[WIDTH*389+:WIDTH]=2.0**16*0.07477164;
k[WIDTH*390+:WIDTH]=2.0**16*-0.02643722;
k[WIDTH*391+:WIDTH]=2.0**16*0.06743621;
k[WIDTH*392+:WIDTH]=2.0**16*0.03446252;
k[WIDTH*393+:WIDTH]=2.0**16*-0.08266958;
k[WIDTH*394+:WIDTH]=2.0**16*0.01596777;
k[WIDTH*395+:WIDTH]=2.0**16*-0.08107528;
k[WIDTH*396+:WIDTH]=2.0**16*0.07438820;
k[WIDTH*397+:WIDTH]=2.0**16*0.09107419;
k[WIDTH*398+:WIDTH]=2.0**16*0.05046712;
k[WIDTH*399+:WIDTH]=2.0**16*0.10214583;
k[WIDTH*400+:WIDTH]=2.0**16*0.05047948;
k[WIDTH*401+:WIDTH]=2.0**16*0.00518114;
k[WIDTH*402+:WIDTH]=2.0**16*-0.07588737;
k[WIDTH*403+:WIDTH]=2.0**16*0.00888282;
k[WIDTH*404+:WIDTH]=2.0**16*-0.02132849;
k[WIDTH*405+:WIDTH]=2.0**16*0.03125162;
k[WIDTH*406+:WIDTH]=2.0**16*-0.00487092;
k[WIDTH*407+:WIDTH]=2.0**16*-0.03602469;
k[WIDTH*408+:WIDTH]=2.0**16*0.00703374;
k[WIDTH*409+:WIDTH]=2.0**16*0.06401423;
k[WIDTH*410+:WIDTH]=2.0**16*0.03853321;
k[WIDTH*411+:WIDTH]=2.0**16*0.03531087;
k[WIDTH*412+:WIDTH]=2.0**16*0.03355344;
k[WIDTH*413+:WIDTH]=2.0**16*0.01364304;
k[WIDTH*414+:WIDTH]=2.0**16*0.02529657;
k[WIDTH*415+:WIDTH]=2.0**16*-0.00241210;
k[WIDTH*416+:WIDTH]=2.0**16*0.01443078;
k[WIDTH*417+:WIDTH]=2.0**16*-0.00419206;
k[WIDTH*418+:WIDTH]=2.0**16*-0.04620698;
k[WIDTH*419+:WIDTH]=2.0**16*0.01902756;
k[WIDTH*420+:WIDTH]=2.0**16*0.09754718;
k[WIDTH*421+:WIDTH]=2.0**16*-0.05222283;
k[WIDTH*422+:WIDTH]=2.0**16*0.11522151;
k[WIDTH*423+:WIDTH]=2.0**16*-0.00422172;
k[WIDTH*424+:WIDTH]=2.0**16*0.02531072;
k[WIDTH*425+:WIDTH]=2.0**16*0.00079438;
k[WIDTH*426+:WIDTH]=2.0**16*0.04277046;
k[WIDTH*427+:WIDTH]=2.0**16*-0.10576923;
k[WIDTH*428+:WIDTH]=2.0**16*0.05815171;
k[WIDTH*429+:WIDTH]=2.0**16*-0.04300173;
k[WIDTH*430+:WIDTH]=2.0**16*-0.00655255;
k[WIDTH*431+:WIDTH]=2.0**16*0.02005037;
k[WIDTH*432+:WIDTH]=2.0**16*-0.04184856;
k[WIDTH*433+:WIDTH]=2.0**16*0.01855580;
k[WIDTH*434+:WIDTH]=2.0**16*0.07405847;
k[WIDTH*435+:WIDTH]=2.0**16*0.02127345;
k[WIDTH*436+:WIDTH]=2.0**16*-0.04189354;
k[WIDTH*437+:WIDTH]=2.0**16*-0.02086769;
k[WIDTH*438+:WIDTH]=2.0**16*-0.09067781;
k[WIDTH*439+:WIDTH]=2.0**16*0.02463831;
k[WIDTH*440+:WIDTH]=2.0**16*0.02951787;
k[WIDTH*441+:WIDTH]=2.0**16*-0.10920864;
k[WIDTH*442+:WIDTH]=2.0**16*0.05734766;
k[WIDTH*443+:WIDTH]=2.0**16*0.02487890;
k[WIDTH*444+:WIDTH]=2.0**16*-0.00051090;
k[WIDTH*445+:WIDTH]=2.0**16*-0.01192762;
k[WIDTH*446+:WIDTH]=2.0**16*0.02244899;
k[WIDTH*447+:WIDTH]=2.0**16*0.18104414;
k[WIDTH*448+:WIDTH]=2.0**16*0.01822764;
k[WIDTH*449+:WIDTH]=2.0**16*-0.03158866;
k[WIDTH*450+:WIDTH]=2.0**16*0.03746881;
k[WIDTH*451+:WIDTH]=2.0**16*0.01583556;
k[WIDTH*452+:WIDTH]=2.0**16*-0.01378931;
k[WIDTH*453+:WIDTH]=2.0**16*0.00157250;
k[WIDTH*454+:WIDTH]=2.0**16*-0.09839753;
k[WIDTH*455+:WIDTH]=2.0**16*0.00396166;
k[WIDTH*456+:WIDTH]=2.0**16*0.01842272;
k[WIDTH*457+:WIDTH]=2.0**16*-0.08265156;
k[WIDTH*458+:WIDTH]=2.0**16*0.04101302;
k[WIDTH*459+:WIDTH]=2.0**16*0.09889290;
k[WIDTH*460+:WIDTH]=2.0**16*-0.01738016;
k[WIDTH*461+:WIDTH]=2.0**16*-0.08669725;
k[WIDTH*462+:WIDTH]=2.0**16*-0.03378740;
k[WIDTH*463+:WIDTH]=2.0**16*-0.01905030;
k[WIDTH*464+:WIDTH]=2.0**16*0.00349438;
k[WIDTH*465+:WIDTH]=2.0**16*-0.02029700;
k[WIDTH*466+:WIDTH]=2.0**16*0.05208898;
k[WIDTH*467+:WIDTH]=2.0**16*-0.03173044;
k[WIDTH*468+:WIDTH]=2.0**16*-0.02375421;
k[WIDTH*469+:WIDTH]=2.0**16*0.01592865;
k[WIDTH*470+:WIDTH]=2.0**16*0.09345986;
k[WIDTH*471+:WIDTH]=2.0**16*0.06100347;
k[WIDTH*472+:WIDTH]=2.0**16*0.05674489;
k[WIDTH*473+:WIDTH]=2.0**16*-0.01168999;
k[WIDTH*474+:WIDTH]=2.0**16*-0.00549902;
k[WIDTH*475+:WIDTH]=2.0**16*-0.03355075;
k[WIDTH*476+:WIDTH]=2.0**16*-0.07697343;
k[WIDTH*477+:WIDTH]=2.0**16*0.07342120;
k[WIDTH*478+:WIDTH]=2.0**16*0.09126708;
k[WIDTH*479+:WIDTH]=2.0**16*-0.06468960;
k[WIDTH*480+:WIDTH]=2.0**16*0.06964764;
k[WIDTH*481+:WIDTH]=2.0**16*0.03985672;
k[WIDTH*482+:WIDTH]=2.0**16*-0.05352214;
k[WIDTH*483+:WIDTH]=2.0**16*-0.01221178;
k[WIDTH*484+:WIDTH]=2.0**16*0.03479894;
k[WIDTH*485+:WIDTH]=2.0**16*-0.02537390;
k[WIDTH*486+:WIDTH]=2.0**16*0.09487378;
k[WIDTH*487+:WIDTH]=2.0**16*-0.03637711;
k[WIDTH*488+:WIDTH]=2.0**16*-0.00922548;
k[WIDTH*489+:WIDTH]=2.0**16*0.10492546;
k[WIDTH*490+:WIDTH]=2.0**16*-0.02407874;
k[WIDTH*491+:WIDTH]=2.0**16*0.06734608;
k[WIDTH*492+:WIDTH]=2.0**16*0.05578750;
k[WIDTH*493+:WIDTH]=2.0**16*-0.03725347;
k[WIDTH*494+:WIDTH]=2.0**16*-0.03501960;
k[WIDTH*495+:WIDTH]=2.0**16*-0.07208083;
k[WIDTH*496+:WIDTH]=2.0**16*-0.01665732;
k[WIDTH*497+:WIDTH]=2.0**16*0.05019510;
k[WIDTH*498+:WIDTH]=2.0**16*-0.00314929;
k[WIDTH*499+:WIDTH]=2.0**16*-0.00345129;
k[WIDTH*500+:WIDTH]=2.0**16*-0.03605704;
k[WIDTH*501+:WIDTH]=2.0**16*0.00286291;
k[WIDTH*502+:WIDTH]=2.0**16*-0.00890034;
k[WIDTH*503+:WIDTH]=2.0**16*-0.03926211;
k[WIDTH*504+:WIDTH]=2.0**16*-0.03774858;
k[WIDTH*505+:WIDTH]=2.0**16*0.04859263;
k[WIDTH*506+:WIDTH]=2.0**16*-0.05835532;
k[WIDTH*507+:WIDTH]=2.0**16*0.02726348;
k[WIDTH*508+:WIDTH]=2.0**16*0.04084381;
k[WIDTH*509+:WIDTH]=2.0**16*0.04991816;
k[WIDTH*510+:WIDTH]=2.0**16*-0.02580752;
k[WIDTH*511+:WIDTH]=2.0**16*-0.03771202;
	end
	endtask
	
	task initb;
	begin
b[WIDTH*0+:WIDTH]=2.0**16*-8.63873340;
b[WIDTH*1+:WIDTH]=2.0**16*-327.04871179;
b[WIDTH*2+:WIDTH]=2.0**16*-64.78867382;
b[WIDTH*3+:WIDTH]=2.0**16*-71.99319358;
b[WIDTH*4+:WIDTH]=2.0**16*80.14839894;
b[WIDTH*5+:WIDTH]=2.0**16*104.41575475;
b[WIDTH*6+:WIDTH]=2.0**16*-56.26097181;
b[WIDTH*7+:WIDTH]=2.0**16*-156.31807115;
b[WIDTH*8+:WIDTH]=2.0**16*-214.47508655;
b[WIDTH*9+:WIDTH]=2.0**16*-4.57304511;
b[WIDTH*10+:WIDTH]=2.0**16*-63.54444655;
b[WIDTH*11+:WIDTH]=2.0**16*-232.06578039;
b[WIDTH*12+:WIDTH]=2.0**16*-38.60679546;
b[WIDTH*13+:WIDTH]=2.0**16*-64.49636815;
b[WIDTH*14+:WIDTH]=2.0**16*-99.12426097;
b[WIDTH*15+:WIDTH]=2.0**16*3.70355178;
b[WIDTH*16+:WIDTH]=2.0**16*135.89150321;
b[WIDTH*17+:WIDTH]=2.0**16*-41.18853471;
b[WIDTH*18+:WIDTH]=2.0**16*-208.64555269;
b[WIDTH*19+:WIDTH]=2.0**16*90.28606468;
b[WIDTH*20+:WIDTH]=2.0**16*-244.30680251;
b[WIDTH*21+:WIDTH]=2.0**16*-19.44543639;
b[WIDTH*22+:WIDTH]=2.0**16*85.54237970;
b[WIDTH*23+:WIDTH]=2.0**16*-13.57849358;
b[WIDTH*24+:WIDTH]=2.0**16*185.14760462;
b[WIDTH*25+:WIDTH]=2.0**16*133.88763289;
b[WIDTH*26+:WIDTH]=2.0**16*-60.43698785;
b[WIDTH*27+:WIDTH]=2.0**16*160.90274458;
b[WIDTH*28+:WIDTH]=2.0**16*-59.76158762;
b[WIDTH*29+:WIDTH]=2.0**16*188.43205337;
b[WIDTH*30+:WIDTH]=2.0**16*24.28932399;
b[WIDTH*31+:WIDTH]=2.0**16*27.74813956;
	end
	endtask
	
	task inita;
	begin
a[WIDTH*0+:WIDTH]=2.0**16*0.53766714;
a[WIDTH*1+:WIDTH]=2.0**16*-1.06887046;
a[WIDTH*2+:WIDTH]=2.0**16*1.54421190;
a[WIDTH*3+:WIDTH]=2.0**16*-0.08249443;
a[WIDTH*4+:WIDTH]=2.0**16*0.70154146;
a[WIDTH*5+:WIDTH]=2.0**16*-0.29375360;
a[WIDTH*6+:WIDTH]=2.0**16*-0.30310762;
a[WIDTH*7+:WIDTH]=2.0**16*-1.50615970;
a[WIDTH*8+:WIDTH]=2.0**16*2.02369089;
a[WIDTH*9+:WIDTH]=2.0**16*1.19210187;
a[WIDTH*10+:WIDTH]=2.0**16*-1.01494364;
a[WIDTH*11+:WIDTH]=2.0**16*-0.78414618;
a[WIDTH*12+:WIDTH]=2.0**16*-1.03598478;
a[WIDTH*13+:WIDTH]=2.0**16*-0.29258813;
a[WIDTH*14+:WIDTH]=2.0**16*-0.42505849;
a[WIDTH*15+:WIDTH]=2.0**16*0.17694682;
a[WIDTH*16+:WIDTH]=2.0**16*1.83388501;
a[WIDTH*17+:WIDTH]=2.0**16*-0.80949869;
a[WIDTH*18+:WIDTH]=2.0**16*0.08593113;
a[WIDTH*19+:WIDTH]=2.0**16*-1.93302292;
a[WIDTH*20+:WIDTH]=2.0**16*-2.05181630;
a[WIDTH*21+:WIDTH]=2.0**16*-0.84792624;
a[WIDTH*22+:WIDTH]=2.0**16*0.02304562;
a[WIDTH*23+:WIDTH]=2.0**16*-0.44462782;
a[WIDTH*24+:WIDTH]=2.0**16*-2.25835397;
a[WIDTH*25+:WIDTH]=2.0**16*-1.61183039;
a[WIDTH*26+:WIDTH]=2.0**16*-0.47106991;
a[WIDTH*27+:WIDTH]=2.0**16*-1.80537335;
a[WIDTH*28+:WIDTH]=2.0**16*1.87786546;
a[WIDTH*29+:WIDTH]=2.0**16*-0.54078642;
a[WIDTH*30+:WIDTH]=2.0**16*0.58943337;
a[WIDTH*31+:WIDTH]=2.0**16*-0.30750347;
a[WIDTH*32+:WIDTH]=2.0**16*-2.25884686;
a[WIDTH*33+:WIDTH]=2.0**16*-2.94428416;
a[WIDTH*34+:WIDTH]=2.0**16*-1.49159031;
a[WIDTH*35+:WIDTH]=2.0**16*-0.43896615;
a[WIDTH*36+:WIDTH]=2.0**16*-0.35385000;
a[WIDTH*37+:WIDTH]=2.0**16*-1.12012830;
a[WIDTH*38+:WIDTH]=2.0**16*0.05129036;
a[WIDTH*39+:WIDTH]=2.0**16*-0.15594104;
a[WIDTH*40+:WIDTH]=2.0**16*2.22944568;
a[WIDTH*41+:WIDTH]=2.0**16*-0.02446194;
a[WIDTH*42+:WIDTH]=2.0**16*0.13702487;
a[WIDTH*43+:WIDTH]=2.0**16*1.85859295;
a[WIDTH*44+:WIDTH]=2.0**16*0.94070440;
a[WIDTH*45+:WIDTH]=2.0**16*-0.30864182;
a[WIDTH*46+:WIDTH]=2.0**16*-0.06279123;
a[WIDTH*47+:WIDTH]=2.0**16*-0.13182035;
a[WIDTH*48+:WIDTH]=2.0**16*0.86217332;
a[WIDTH*49+:WIDTH]=2.0**16*1.43838029;
a[WIDTH*50+:WIDTH]=2.0**16*-0.74230184;
a[WIDTH*51+:WIDTH]=2.0**16*-1.79467884;
a[WIDTH*52+:WIDTH]=2.0**16*-0.82358653;
a[WIDTH*53+:WIDTH]=2.0**16*2.52599969;
a[WIDTH*54+:WIDTH]=2.0**16*0.82606279;
a[WIDTH*55+:WIDTH]=2.0**16*0.27606825;
a[WIDTH*56+:WIDTH]=2.0**16*0.33756370;
a[WIDTH*57+:WIDTH]=2.0**16*-1.94884718;
a[WIDTH*58+:WIDTH]=2.0**16*-0.29186338;
a[WIDTH*59+:WIDTH]=2.0**16*-0.60453009;
a[WIDTH*60+:WIDTH]=2.0**16*0.78734578;
a[WIDTH*61+:WIDTH]=2.0**16*-1.09659330;
a[WIDTH*62+:WIDTH]=2.0**16*-2.02195893;
a[WIDTH*63+:WIDTH]=2.0**16*0.59535767;
a[WIDTH*64+:WIDTH]=2.0**16*0.31876524;
a[WIDTH*65+:WIDTH]=2.0**16*0.32519054;
a[WIDTH*66+:WIDTH]=2.0**16*-1.06158173;
a[WIDTH*67+:WIDTH]=2.0**16*0.84037553;
a[WIDTH*68+:WIDTH]=2.0**16*-1.57705702;
a[WIDTH*69+:WIDTH]=2.0**16*1.65549759;
a[WIDTH*70+:WIDTH]=2.0**16*1.52697669;
a[WIDTH*71+:WIDTH]=2.0**16*-0.26116365;
a[WIDTH*72+:WIDTH]=2.0**16*1.00006082;
a[WIDTH*73+:WIDTH]=2.0**16*1.02049801;
a[WIDTH*74+:WIDTH]=2.0**16*0.30181856;
a[WIDTH*75+:WIDTH]=2.0**16*0.10335972;
a[WIDTH*76+:WIDTH]=2.0**16*-0.87587426;
a[WIDTH*77+:WIDTH]=2.0**16*-0.49300982;
a[WIDTH*78+:WIDTH]=2.0**16*-0.98213153;
a[WIDTH*79+:WIDTH]=2.0**16*1.04683278;
a[WIDTH*80+:WIDTH]=2.0**16*-1.30768830;
a[WIDTH*81+:WIDTH]=2.0**16*-0.75492832;
a[WIDTH*82+:WIDTH]=2.0**16*2.35045722;
a[WIDTH*83+:WIDTH]=2.0**16*-0.88803208;
a[WIDTH*84+:WIDTH]=2.0**16*0.50797465;
a[WIDTH*85+:WIDTH]=2.0**16*0.30753516;
a[WIDTH*86+:WIDTH]=2.0**16*0.46691444;
a[WIDTH*87+:WIDTH]=2.0**16*0.44342191;
a[WIDTH*88+:WIDTH]=2.0**16*-1.66416447;
a[WIDTH*89+:WIDTH]=2.0**16*0.86171630;
a[WIDTH*90+:WIDTH]=2.0**16*0.39993094;
a[WIDTH*91+:WIDTH]=2.0**16*0.56316696;
a[WIDTH*92+:WIDTH]=2.0**16*0.31994913;
a[WIDTH*93+:WIDTH]=2.0**16*-0.18073936;
a[WIDTH*94+:WIDTH]=2.0**16*0.61251130;
a[WIDTH*95+:WIDTH]=2.0**16*-0.19795863;
a[WIDTH*96+:WIDTH]=2.0**16*-0.43359202;
a[WIDTH*97+:WIDTH]=2.0**16*1.37029854;
a[WIDTH*98+:WIDTH]=2.0**16*-0.61560188;
a[WIDTH*99+:WIDTH]=2.0**16*0.10009283;
a[WIDTH*100+:WIDTH]=2.0**16*0.28198406;
a[WIDTH*101+:WIDTH]=2.0**16*-1.25711836;
a[WIDTH*102+:WIDTH]=2.0**16*-0.20971334;
a[WIDTH*103+:WIDTH]=2.0**16*0.39189421;
a[WIDTH*104+:WIDTH]=2.0**16*-0.59003456;
a[WIDTH*105+:WIDTH]=2.0**16*0.00116208;
a[WIDTH*106+:WIDTH]=2.0**16*-0.92996156;
a[WIDTH*107+:WIDTH]=2.0**16*0.11359700;
a[WIDTH*108+:WIDTH]=2.0**16*-0.55829428;
a[WIDTH*109+:WIDTH]=2.0**16*0.04584111;
a[WIDTH*110+:WIDTH]=2.0**16*-0.05488613;
a[WIDTH*111+:WIDTH]=2.0**16*0.32767816;
a[WIDTH*112+:WIDTH]=2.0**16*0.34262447;
a[WIDTH*113+:WIDTH]=2.0**16*-1.71151642;
a[WIDTH*114+:WIDTH]=2.0**16*0.74807678;
a[WIDTH*115+:WIDTH]=2.0**16*-0.54452893;
a[WIDTH*116+:WIDTH]=2.0**16*0.03347988;
a[WIDTH*117+:WIDTH]=2.0**16*-0.86546803;
a[WIDTH*118+:WIDTH]=2.0**16*0.62519036;
a[WIDTH*119+:WIDTH]=2.0**16*-1.25067891;
a[WIDTH*120+:WIDTH]=2.0**16*-0.27806416;
a[WIDTH*121+:WIDTH]=2.0**16*-0.07083721;
a[WIDTH*122+:WIDTH]=2.0**16*-0.17683027;
a[WIDTH*123+:WIDTH]=2.0**16*-0.90472621;
a[WIDTH*124+:WIDTH]=2.0**16*-0.31142942;
a[WIDTH*125+:WIDTH]=2.0**16*-0.06378312;
a[WIDTH*126+:WIDTH]=2.0**16*-1.11873200;
a[WIDTH*127+:WIDTH]=2.0**16*-0.23830150;
a[WIDTH*128+:WIDTH]=2.0**16*3.57839694;
a[WIDTH*129+:WIDTH]=2.0**16*-0.10224245;
a[WIDTH*130+:WIDTH]=2.0**16*-0.19241851;
a[WIDTH*131+:WIDTH]=2.0**16*0.30352079;
a[WIDTH*132+:WIDTH]=2.0**16*-1.33367794;
a[WIDTH*133+:WIDTH]=2.0**16*-0.17653411;
a[WIDTH*134+:WIDTH]=2.0**16*0.18322726;
a[WIDTH*135+:WIDTH]=2.0**16*-0.94796092;
a[WIDTH*136+:WIDTH]=2.0**16*0.42271569;
a[WIDTH*137+:WIDTH]=2.0**16*-2.48628392;
a[WIDTH*138+:WIDTH]=2.0**16*-2.13209460;
a[WIDTH*139+:WIDTH]=2.0**16*-0.46771458;
a[WIDTH*140+:WIDTH]=2.0**16*-0.57000992;
a[WIDTH*141+:WIDTH]=2.0**16*0.61133519;
a[WIDTH*142+:WIDTH]=2.0**16*-0.62637854;
a[WIDTH*143+:WIDTH]=2.0**16*0.22959689;
a[WIDTH*144+:WIDTH]=2.0**16*2.76943703;
a[WIDTH*145+:WIDTH]=2.0**16*-0.24144704;
a[WIDTH*146+:WIDTH]=2.0**16*0.88861043;
a[WIDTH*147+:WIDTH]=2.0**16*-0.60032656;
a[WIDTH*148+:WIDTH]=2.0**16*1.12749228;
a[WIDTH*149+:WIDTH]=2.0**16*0.79141606;
a[WIDTH*150+:WIDTH]=2.0**16*-1.02976754;
a[WIDTH*151+:WIDTH]=2.0**16*-0.74110609;
a[WIDTH*152+:WIDTH]=2.0**16*-1.67020070;
a[WIDTH*153+:WIDTH]=2.0**16*0.58117232;
a[WIDTH*154+:WIDTH]=2.0**16*1.14536171;
a[WIDTH*155+:WIDTH]=2.0**16*-0.12488995;
a[WIDTH*156+:WIDTH]=2.0**16*-1.02573362;
a[WIDTH*157+:WIDTH]=2.0**16*0.10931769;
a[WIDTH*158+:WIDTH]=2.0**16*0.24951774;
a[WIDTH*159+:WIDTH]=2.0**16*0.43999790;
a[WIDTH*160+:WIDTH]=2.0**16*-1.34988694;
a[WIDTH*161+:WIDTH]=2.0**16*0.31920674;
a[WIDTH*162+:WIDTH]=2.0**16*-0.76484924;
a[WIDTH*163+:WIDTH]=2.0**16*0.48996532;
a[WIDTH*164+:WIDTH]=2.0**16*0.35017941;
a[WIDTH*165+:WIDTH]=2.0**16*-1.33200442;
a[WIDTH*166+:WIDTH]=2.0**16*0.94922183;
a[WIDTH*167+:WIDTH]=2.0**16*-0.50781755;
a[WIDTH*168+:WIDTH]=2.0**16*0.47163433;
a[WIDTH*169+:WIDTH]=2.0**16*-2.19243492;
a[WIDTH*170+:WIDTH]=2.0**16*-0.62909076;
a[WIDTH*171+:WIDTH]=2.0**16*1.47895849;
a[WIDTH*172+:WIDTH]=2.0**16*-0.90874559;
a[WIDTH*173+:WIDTH]=2.0**16*1.81401545;
a[WIDTH*174+:WIDTH]=2.0**16*-0.99301901;
a[WIDTH*175+:WIDTH]=2.0**16*-0.61686593;
a[WIDTH*176+:WIDTH]=2.0**16*3.03492347;
a[WIDTH*177+:WIDTH]=2.0**16*0.31285860;
a[WIDTH*178+:WIDTH]=2.0**16*-1.40226897;
a[WIDTH*179+:WIDTH]=2.0**16*0.73936312;
a[WIDTH*180+:WIDTH]=2.0**16*-0.29906603;
a[WIDTH*181+:WIDTH]=2.0**16*-2.32986716;
a[WIDTH*182+:WIDTH]=2.0**16*0.30706192;
a[WIDTH*183+:WIDTH]=2.0**16*-0.32057551;
a[WIDTH*184+:WIDTH]=2.0**16*-1.21284720;
a[WIDTH*185+:WIDTH]=2.0**16*-2.31928031;
a[WIDTH*186+:WIDTH]=2.0**16*-1.20384997;
a[WIDTH*187+:WIDTH]=2.0**16*-0.86081569;
a[WIDTH*188+:WIDTH]=2.0**16*-0.20989733;
a[WIDTH*189+:WIDTH]=2.0**16*0.31202383;
a[WIDTH*190+:WIDTH]=2.0**16*0.97495022;
a[WIDTH*191+:WIDTH]=2.0**16*0.27483679;
a[WIDTH*192+:WIDTH]=2.0**16*0.72540422;
a[WIDTH*193+:WIDTH]=2.0**16*-0.86487992;
a[WIDTH*194+:WIDTH]=2.0**16*-1.42237593;
a[WIDTH*195+:WIDTH]=2.0**16*1.71188778;
a[WIDTH*196+:WIDTH]=2.0**16*0.02288979;
a[WIDTH*197+:WIDTH]=2.0**16*-1.44909729;
a[WIDTH*198+:WIDTH]=2.0**16*0.13517494;
a[WIDTH*199+:WIDTH]=2.0**16*0.01246904;
a[WIDTH*200+:WIDTH]=2.0**16*0.06619005;
a[WIDTH*201+:WIDTH]=2.0**16*0.07993371;
a[WIDTH*202+:WIDTH]=2.0**16*-0.25394468;
a[WIDTH*203+:WIDTH]=2.0**16*0.78466847;
a[WIDTH*204+:WIDTH]=2.0**16*-1.69886408;
a[WIDTH*205+:WIDTH]=2.0**16*1.80449377;
a[WIDTH*206+:WIDTH]=2.0**16*-0.64070951;
a[WIDTH*207+:WIDTH]=2.0**16*0.60110203;
a[WIDTH*208+:WIDTH]=2.0**16*-0.06305487;
a[WIDTH*209+:WIDTH]=2.0**16*-0.03005130;
a[WIDTH*210+:WIDTH]=2.0**16*0.48819391;
a[WIDTH*211+:WIDTH]=2.0**16*-0.19412354;
a[WIDTH*212+:WIDTH]=2.0**16*-0.26199543;
a[WIDTH*213+:WIDTH]=2.0**16*0.33351083;
a[WIDTH*214+:WIDTH]=2.0**16*0.51524634;
a[WIDTH*215+:WIDTH]=2.0**16*-3.02917734;
a[WIDTH*216+:WIDTH]=2.0**16*0.65235589;
a[WIDTH*217+:WIDTH]=2.0**16*-0.94848098;
a[WIDTH*218+:WIDTH]=2.0**16*-1.42864686;
a[WIDTH*219+:WIDTH]=2.0**16*0.30862314;
a[WIDTH*220+:WIDTH]=2.0**16*0.60760058;
a[WIDTH*221+:WIDTH]=2.0**16*-0.72312148;
a[WIDTH*222+:WIDTH]=2.0**16*1.80886262;
a[WIDTH*223+:WIDTH]=2.0**16*0.09230795;
a[WIDTH*224+:WIDTH]=2.0**16*0.71474290;
a[WIDTH*225+:WIDTH]=2.0**16*-0.16487902;
a[WIDTH*226+:WIDTH]=2.0**16*-0.17737516;
a[WIDTH*227+:WIDTH]=2.0**16*-2.13835527;
a[WIDTH*228+:WIDTH]=2.0**16*-1.75021237;
a[WIDTH*229+:WIDTH]=2.0**16*0.39135360;
a[WIDTH*230+:WIDTH]=2.0**16*0.26140632;
a[WIDTH*231+:WIDTH]=2.0**16*-0.45701464;
a[WIDTH*232+:WIDTH]=2.0**16*0.32705997;
a[WIDTH*233+:WIDTH]=2.0**16*0.41149062;
a[WIDTH*234+:WIDTH]=2.0**16*-0.02085762;
a[WIDTH*235+:WIDTH]=2.0**16*-0.23386004;
a[WIDTH*236+:WIDTH]=2.0**16*-0.11779829;
a[WIDTH*237+:WIDTH]=2.0**16*0.52654704;
a[WIDTH*238+:WIDTH]=2.0**16*-1.07986625;
a[WIDTH*239+:WIDTH]=2.0**16*1.72984139;
a[WIDTH*240+:WIDTH]=2.0**16*-0.20496606;
a[WIDTH*241+:WIDTH]=2.0**16*0.62770729;
a[WIDTH*242+:WIDTH]=2.0**16*-0.19605349;
a[WIDTH*243+:WIDTH]=2.0**16*-0.83958875;
a[WIDTH*244+:WIDTH]=2.0**16*-0.28565097;
a[WIDTH*245+:WIDTH]=2.0**16*0.45167942;
a[WIDTH*246+:WIDTH]=2.0**16*-0.94148577;
a[WIDTH*247+:WIDTH]=2.0**16*1.24244841;
a[WIDTH*248+:WIDTH]=2.0**16*1.08263350;
a[WIDTH*249+:WIDTH]=2.0**16*0.67697781;
a[WIDTH*250+:WIDTH]=2.0**16*-0.56066500;
a[WIDTH*251+:WIDTH]=2.0**16*-1.05697275;
a[WIDTH*252+:WIDTH]=2.0**16*0.69916033;
a[WIDTH*253+:WIDTH]=2.0**16*-0.26025086;
a[WIDTH*254+:WIDTH]=2.0**16*0.19918944;
a[WIDTH*255+:WIDTH]=2.0**16*-0.60855744;
a[WIDTH*256+:WIDTH]=2.0**16*-0.12414435;
a[WIDTH*257+:WIDTH]=2.0**16*1.09326567;
a[WIDTH*258+:WIDTH]=2.0**16*1.41931015;
a[WIDTH*259+:WIDTH]=2.0**16*1.35459433;
a[WIDTH*260+:WIDTH]=2.0**16*-0.83136651;
a[WIDTH*261+:WIDTH]=2.0**16*-0.13028465;
a[WIDTH*262+:WIDTH]=2.0**16*-0.16233767;
a[WIDTH*263+:WIDTH]=2.0**16*-1.06670140;
a[WIDTH*264+:WIDTH]=2.0**16*1.00607711;
a[WIDTH*265+:WIDTH]=2.0**16*0.85773255;
a[WIDTH*266+:WIDTH]=2.0**16*2.17777871;
a[WIDTH*267+:WIDTH]=2.0**16*-0.28414095;
a[WIDTH*268+:WIDTH]=2.0**16*0.26964864;
a[WIDTH*269+:WIDTH]=2.0**16*0.60014251;
a[WIDTH*270+:WIDTH]=2.0**16*-1.52102656;
a[WIDTH*271+:WIDTH]=2.0**16*-0.73705977;
a[WIDTH*272+:WIDTH]=2.0**16*1.48969761;
a[WIDTH*273+:WIDTH]=2.0**16*1.10927330;
a[WIDTH*274+:WIDTH]=2.0**16*0.29158437;
a[WIDTH*275+:WIDTH]=2.0**16*-1.07215529;
a[WIDTH*276+:WIDTH]=2.0**16*-0.97920631;
a[WIDTH*277+:WIDTH]=2.0**16*0.18368910;
a[WIDTH*278+:WIDTH]=2.0**16*-0.14605463;
a[WIDTH*279+:WIDTH]=2.0**16*0.93372816;
a[WIDTH*280+:WIDTH]=2.0**16*-0.65090774;
a[WIDTH*281+:WIDTH]=2.0**16*-0.69115913;
a[WIDTH*282+:WIDTH]=2.0**16*1.13846539;
a[WIDTH*283+:WIDTH]=2.0**16*-0.08669028;
a[WIDTH*284+:WIDTH]=2.0**16*0.49428706;
a[WIDTH*285+:WIDTH]=2.0**16*0.59393080;
a[WIDTH*286+:WIDTH]=2.0**16*-0.72363113;
a[WIDTH*287+:WIDTH]=2.0**16*-1.74987931;
a[WIDTH*288+:WIDTH]=2.0**16*1.40903449;
a[WIDTH*289+:WIDTH]=2.0**16*-0.86365282;
a[WIDTH*290+:WIDTH]=2.0**16*0.19781105;
a[WIDTH*291+:WIDTH]=2.0**16*0.96095387;
a[WIDTH*292+:WIDTH]=2.0**16*-1.15640166;
a[WIDTH*293+:WIDTH]=2.0**16*-0.47615302;
a[WIDTH*294+:WIDTH]=2.0**16*-0.53201138;
a[WIDTH*295+:WIDTH]=2.0**16*0.35032100;
a[WIDTH*296+:WIDTH]=2.0**16*0.25705616;
a[WIDTH*297+:WIDTH]=2.0**16*0.44937762;
a[WIDTH*298+:WIDTH]=2.0**16*-2.49688650;
a[WIDTH*299+:WIDTH]=2.0**16*-1.46939507;
a[WIDTH*300+:WIDTH]=2.0**16*-1.48312102;
a[WIDTH*301+:WIDTH]=2.0**16*-2.18602161;
a[WIDTH*302+:WIDTH]=2.0**16*-0.59325032;
a[WIDTH*303+:WIDTH]=2.0**16*0.91048258;
a[WIDTH*304+:WIDTH]=2.0**16*1.41719241;
a[WIDTH*305+:WIDTH]=2.0**16*0.07735909;
a[WIDTH*306+:WIDTH]=2.0**16*1.58769909;
a[WIDTH*307+:WIDTH]=2.0**16*0.12404980;
a[WIDTH*308+:WIDTH]=2.0**16*-0.53355711;
a[WIDTH*309+:WIDTH]=2.0**16*0.86202161;
a[WIDTH*310+:WIDTH]=2.0**16*1.68210359;
a[WIDTH*311+:WIDTH]=2.0**16*-0.02900576;
a[WIDTH*312+:WIDTH]=2.0**16*-0.94437781;
a[WIDTH*313+:WIDTH]=2.0**16*0.10063335;
a[WIDTH*314+:WIDTH]=2.0**16*0.44132693;
a[WIDTH*315+:WIDTH]=2.0**16*0.19218224;
a[WIDTH*316+:WIDTH]=2.0**16*-1.02026439;
a[WIDTH*317+:WIDTH]=2.0**16*-1.32704315;
a[WIDTH*318+:WIDTH]=2.0**16*0.40133634;
a[WIDTH*319+:WIDTH]=2.0**16*0.86708255;
a[WIDTH*320+:WIDTH]=2.0**16*0.67149713;
a[WIDTH*321+:WIDTH]=2.0**16*-1.21411704;
a[WIDTH*322+:WIDTH]=2.0**16*-0.80446596;
a[WIDTH*323+:WIDTH]=2.0**16*1.43669662;
a[WIDTH*324+:WIDTH]=2.0**16*-2.00263574;
a[WIDTH*325+:WIDTH]=2.0**16*-1.36169447;
a[WIDTH*326+:WIDTH]=2.0**16*-0.87572935;
a[WIDTH*327+:WIDTH]=2.0**16*0.18245217;
a[WIDTH*328+:WIDTH]=2.0**16*-1.32178852;
a[WIDTH*329+:WIDTH]=2.0**16*0.82607000;
a[WIDTH*330+:WIDTH]=2.0**16*-1.39813788;
a[WIDTH*331+:WIDTH]=2.0**16*-0.82229328;
a[WIDTH*332+:WIDTH]=2.0**16*-0.44699501;
a[WIDTH*333+:WIDTH]=2.0**16*-1.44101360;
a[WIDTH*334+:WIDTH]=2.0**16*0.94213332;
a[WIDTH*335+:WIDTH]=2.0**16*-0.07989284;
a[WIDTH*336+:WIDTH]=2.0**16*-1.20748692;
a[WIDTH*337+:WIDTH]=2.0**16*-1.11350074;
a[WIDTH*338+:WIDTH]=2.0**16*0.69662442;
a[WIDTH*339+:WIDTH]=2.0**16*-1.96090000;
a[WIDTH*340+:WIDTH]=2.0**16*0.96422942;
a[WIDTH*341+:WIDTH]=2.0**16*0.45502956;
a[WIDTH*342+:WIDTH]=2.0**16*-0.48381505;
a[WIDTH*343+:WIDTH]=2.0**16*-1.56505601;
a[WIDTH*344+:WIDTH]=2.0**16*0.92482593;
a[WIDTH*345+:WIDTH]=2.0**16*0.53615708;
a[WIDTH*346+:WIDTH]=2.0**16*-0.25505518;
a[WIDTH*347+:WIDTH]=2.0**16*-0.09424059;
a[WIDTH*348+:WIDTH]=2.0**16*0.10965859;
a[WIDTH*349+:WIDTH]=2.0**16*0.40184450;
a[WIDTH*350+:WIDTH]=2.0**16*0.30048597;
a[WIDTH*351+:WIDTH]=2.0**16*0.89847599;
a[WIDTH*352+:WIDTH]=2.0**16*0.71723865;
a[WIDTH*353+:WIDTH]=2.0**16*-0.00684933;
a[WIDTH*354+:WIDTH]=2.0**16*0.83508817;
a[WIDTH*355+:WIDTH]=2.0**16*-0.19769823;
a[WIDTH*356+:WIDTH]=2.0**16*0.52006010;
a[WIDTH*357+:WIDTH]=2.0**16*-0.84870938;
a[WIDTH*358+:WIDTH]=2.0**16*-0.71200455;
a[WIDTH*359+:WIDTH]=2.0**16*-0.08453948;
a[WIDTH*360+:WIDTH]=2.0**16*0.00004985;
a[WIDTH*361+:WIDTH]=2.0**16*0.89788843;
a[WIDTH*362+:WIDTH]=2.0**16*0.16440407;
a[WIDTH*363+:WIDTH]=2.0**16*0.33621334;
a[WIDTH*364+:WIDTH]=2.0**16*1.12873645;
a[WIDTH*365+:WIDTH]=2.0**16*1.47020128;
a[WIDTH*366+:WIDTH]=2.0**16*-0.37307066;
a[WIDTH*367+:WIDTH]=2.0**16*0.18370342;
a[WIDTH*368+:WIDTH]=2.0**16*1.63023529;
a[WIDTH*369+:WIDTH]=2.0**16*1.53263031;
a[WIDTH*370+:WIDTH]=2.0**16*-0.24371514;
a[WIDTH*371+:WIDTH]=2.0**16*-1.20784549;
a[WIDTH*372+:WIDTH]=2.0**16*-0.02002785;
a[WIDTH*373+:WIDTH]=2.0**16*-0.33488694;
a[WIDTH*374+:WIDTH]=2.0**16*-1.17421233;
a[WIDTH*375+:WIDTH]=2.0**16*1.60394635;
a[WIDTH*376+:WIDTH]=2.0**16*-0.05491891;
a[WIDTH*377+:WIDTH]=2.0**16*-0.13193787;
a[WIDTH*378+:WIDTH]=2.0**16*0.74773403;
a[WIDTH*379+:WIDTH]=2.0**16*-0.90465406;
a[WIDTH*380+:WIDTH]=2.0**16*-0.28996304;
a[WIDTH*381+:WIDTH]=2.0**16*-0.32681423;
a[WIDTH*382+:WIDTH]=2.0**16*0.81548851;
a[WIDTH*383+:WIDTH]=2.0**16*0.29079013;
a[WIDTH*384+:WIDTH]=2.0**16*0.48889377;
a[WIDTH*385+:WIDTH]=2.0**16*-0.76966591;
a[WIDTH*386+:WIDTH]=2.0**16*0.21567009;
a[WIDTH*387+:WIDTH]=2.0**16*2.90800803;
a[WIDTH*388+:WIDTH]=2.0**16*-0.03477109;
a[WIDTH*389+:WIDTH]=2.0**16*0.55278335;
a[WIDTH*390+:WIDTH]=2.0**16*-0.19223952;
a[WIDTH*391+:WIDTH]=2.0**16*0.09834777;
a[WIDTH*392+:WIDTH]=2.0**16*0.91112727;
a[WIDTH*393+:WIDTH]=2.0**16*-0.14720146;
a[WIDTH*394+:WIDTH]=2.0**16*-0.27304695;
a[WIDTH*395+:WIDTH]=2.0**16*-0.28825636;
a[WIDTH*396+:WIDTH]=2.0**16*1.26155072;
a[WIDTH*397+:WIDTH]=2.0**16*0.81232300;
a[WIDTH*398+:WIDTH]=2.0**16*0.79888699;
a[WIDTH*399+:WIDTH]=2.0**16*0.11294472;
a[WIDTH*400+:WIDTH]=2.0**16*1.03469301;
a[WIDTH*401+:WIDTH]=2.0**16*0.37137881;
a[WIDTH*402+:WIDTH]=2.0**16*-1.16584393;
a[WIDTH*403+:WIDTH]=2.0**16*0.82521889;
a[WIDTH*404+:WIDTH]=2.0**16*-0.79816358;
a[WIDTH*405+:WIDTH]=2.0**16*1.03909065;
a[WIDTH*406+:WIDTH]=2.0**16*-0.27407023;
a[WIDTH*407+:WIDTH]=2.0**16*0.04137361;
a[WIDTH*408+:WIDTH]=2.0**16*0.59458370;
a[WIDTH*409+:WIDTH]=2.0**16*1.00777341;
a[WIDTH*410+:WIDTH]=2.0**16*1.57630015;
a[WIDTH*411+:WIDTH]=2.0**16*0.35006276;
a[WIDTH*412+:WIDTH]=2.0**16*0.47542481;
a[WIDTH*413+:WIDTH]=2.0**16*0.54554010;
a[WIDTH*414+:WIDTH]=2.0**16*0.12020528;
a[WIDTH*415+:WIDTH]=2.0**16*0.43995219;
a[WIDTH*416+:WIDTH]=2.0**16*0.72688513;
a[WIDTH*417+:WIDTH]=2.0**16*-0.22558440;
a[WIDTH*418+:WIDTH]=2.0**16*-1.14795278;
a[WIDTH*419+:WIDTH]=2.0**16*1.37897198;
a[WIDTH*420+:WIDTH]=2.0**16*1.01868528;
a[WIDTH*421+:WIDTH]=2.0**16*-1.11763868;
a[WIDTH*422+:WIDTH]=2.0**16*1.53007251;
a[WIDTH*423+:WIDTH]=2.0**16*-0.73416911;
a[WIDTH*424+:WIDTH]=2.0**16*0.35020117;
a[WIDTH*425+:WIDTH]=2.0**16*-2.12365546;
a[WIDTH*426+:WIDTH]=2.0**16*-0.48093715;
a[WIDTH*427+:WIDTH]=2.0**16*-1.83585914;
a[WIDTH*428+:WIDTH]=2.0**16*1.17411675;
a[WIDTH*429+:WIDTH]=2.0**16*-1.05163231;
a[WIDTH*430+:WIDTH]=2.0**16*0.57124763;
a[WIDTH*431+:WIDTH]=2.0**16*0.10166244;
a[WIDTH*432+:WIDTH]=2.0**16*-0.30344092;
a[WIDTH*433+:WIDTH]=2.0**16*1.11735614;
a[WIDTH*434+:WIDTH]=2.0**16*0.10487472;
a[WIDTH*435+:WIDTH]=2.0**16*-1.05818026;
a[WIDTH*436+:WIDTH]=2.0**16*-0.13321748;
a[WIDTH*437+:WIDTH]=2.0**16*1.26065871;
a[WIDTH*438+:WIDTH]=2.0**16*-0.24902474;
a[WIDTH*439+:WIDTH]=2.0**16*-0.03081373;
a[WIDTH*440+:WIDTH]=2.0**16*1.25025123;
a[WIDTH*441+:WIDTH]=2.0**16*-0.50458641;
a[WIDTH*442+:WIDTH]=2.0**16*0.32751212;
a[WIDTH*443+:WIDTH]=2.0**16*1.03597591;
a[WIDTH*444+:WIDTH]=2.0**16*0.12694707;
a[WIDTH*445+:WIDTH]=2.0**16*0.39746700;
a[WIDTH*446+:WIDTH]=2.0**16*0.41279601;
a[WIDTH*447+:WIDTH]=2.0**16*2.78733523;
a[WIDTH*448+:WIDTH]=2.0**16*0.29387147;
a[WIDTH*449+:WIDTH]=2.0**16*-1.08906430;
a[WIDTH*450+:WIDTH]=2.0**16*0.72225403;
a[WIDTH*451+:WIDTH]=2.0**16*-0.46861558;
a[WIDTH*452+:WIDTH]=2.0**16*-0.71453016;
a[WIDTH*453+:WIDTH]=2.0**16*0.66014314;
a[WIDTH*454+:WIDTH]=2.0**16*-1.06421341;
a[WIDTH*455+:WIDTH]=2.0**16*0.23234701;
a[WIDTH*456+:WIDTH]=2.0**16*0.92978946;
a[WIDTH*457+:WIDTH]=2.0**16*-1.27059445;
a[WIDTH*458+:WIDTH]=2.0**16*0.66473412;
a[WIDTH*459+:WIDTH]=2.0**16*2.42446114;
a[WIDTH*460+:WIDTH]=2.0**16*-0.65681593;
a[WIDTH*461+:WIDTH]=2.0**16*-0.75189474;
a[WIDTH*462+:WIDTH]=2.0**16*-0.98696188;
a[WIDTH*463+:WIDTH]=2.0**16*-1.16666503;
a[WIDTH*464+:WIDTH]=2.0**16*-0.78728280;
a[WIDTH*465+:WIDTH]=2.0**16*0.03255746;
a[WIDTH*466+:WIDTH]=2.0**16*2.58549125;
a[WIDTH*467+:WIDTH]=2.0**16*-0.27246941;
a[WIDTH*468+:WIDTH]=2.0**16*1.35138577;
a[WIDTH*469+:WIDTH]=2.0**16*-0.06786555;
a[WIDTH*470+:WIDTH]=2.0**16*1.60345730;
a[WIDTH*471+:WIDTH]=2.0**16*0.42638756;
a[WIDTH*472+:WIDTH]=2.0**16*0.23976326;
a[WIDTH*473+:WIDTH]=2.0**16*-0.38258480;
a[WIDTH*474+:WIDTH]=2.0**16*0.08518859;
a[WIDTH*475+:WIDTH]=2.0**16*0.95940051;
a[WIDTH*476+:WIDTH]=2.0**16*-1.48139907;
a[WIDTH*477+:WIDTH]=2.0**16*1.51626690;
a[WIDTH*478+:WIDTH]=2.0**16*0.75956833;
a[WIDTH*479+:WIDTH]=2.0**16*-1.85429908;
a[WIDTH*480+:WIDTH]=2.0**16*0.88839563;
a[WIDTH*481+:WIDTH]=2.0**16*0.55252702;
a[WIDTH*482+:WIDTH]=2.0**16*-0.66689067;
a[WIDTH*483+:WIDTH]=2.0**16*1.09842462;
a[WIDTH*484+:WIDTH]=2.0**16*-0.22477106;
a[WIDTH*485+:WIDTH]=2.0**16*-0.19522120;
a[WIDTH*486+:WIDTH]=2.0**16*1.23467915;
a[WIDTH*487+:WIDTH]=2.0**16*-0.37280874;
a[WIDTH*488+:WIDTH]=2.0**16*-0.69036110;
a[WIDTH*489+:WIDTH]=2.0**16*0.64867926;
a[WIDTH*490+:WIDTH]=2.0**16*0.88095279;
a[WIDTH*491+:WIDTH]=2.0**16*-0.31577200;
a[WIDTH*492+:WIDTH]=2.0**16*0.15548900;
a[WIDTH*493+:WIDTH]=2.0**16*-0.03256651;
a[WIDTH*494+:WIDTH]=2.0**16*-0.65720130;
a[WIDTH*495+:WIDTH]=2.0**16*-1.14068114;
a[WIDTH*496+:WIDTH]=2.0**16*-1.14707011;
a[WIDTH*497+:WIDTH]=2.0**16*1.10061022;
a[WIDTH*498+:WIDTH]=2.0**16*0.18733102;
a[WIDTH*499+:WIDTH]=2.0**16*-0.27787193;
a[WIDTH*500+:WIDTH]=2.0**16*-0.58902903;
a[WIDTH*501+:WIDTH]=2.0**16*-0.21760635;
a[WIDTH*502+:WIDTH]=2.0**16*-0.22962645;
a[WIDTH*503+:WIDTH]=2.0**16*-0.23645458;
a[WIDTH*504+:WIDTH]=2.0**16*-0.65155364;
a[WIDTH*505+:WIDTH]=2.0**16*0.82572715;
a[WIDTH*506+:WIDTH]=2.0**16*0.32321314;
a[WIDTH*507+:WIDTH]=2.0**16*0.42862268;
a[WIDTH*508+:WIDTH]=2.0**16*0.81855137;
a[WIDTH*509+:WIDTH]=2.0**16*1.63599966;
a[WIDTH*510+:WIDTH]=2.0**16*-0.60391848;
a[WIDTH*511+:WIDTH]=2.0**16*-1.09334346;
	end
	endtask
	
	integer z =0;
	task initx0;
		begin
			for(z=1; z<SIZE; z=z+1) begin
				x0[WIDTH*(SIZE-z)+:WIDTH] = 2**16*1;
			end
			z=1;
		end	
	endtask

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
		x0 = 0;
		k = 0;
		b = 0;
		a = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		$display("START::TiME= ", $time);
		initk;
		inita;
		initb;
		initx0;
		@(posedge clk)
		reset <=1;
		@(posedge clk)
		reset<=0;
		repeat(30*304) begin// 100 clk cycles
			@(posedge clk)
			if(ready) begin
				$display("DONE::TiME= ", $time);
			end
		end
	end
      
endmodule

